`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Last Edits: Nirmal Kumbhare, Ali Akoglu
// 
// Module - data_memory.v
// Description - 32-Bit wide data memory.
//
// INPUTS:-
// Address: 32-Bit address input port.
// WriteData: 32-Bit input port.
// Clk: 1-Bit Input clock signal.
// MemWrite: 1-Bit control signal for memory write.
// MemRead: 1-Bit control signal for memory read.
//
// OUTPUTS:-
// ReadData: 32-Bit registered output port.
//
// FUNCTIONALITY:-
// Design the above memory similar to the 'RegisterFile' model in the previous 
// assignment.  Create a 1K (x32) memory, for which we need 10 bits for the address.  
// In order to implement byte addressing, we will use bits Address[11:2] to index the 
// memory location. 
// The 'WriteData' value is written into the location whose address 
// corresponds to Address[11:2] in the positive clock edge if 'MemWrite' 
// signal is 1. 
// 'ReadData' is the value of memory location Address[11:2] if 
// 'MemRead' is 1, otherwise, it is 0x00000000. The reading of memory is NOT clocked.
//
// you need to declare a 2d array. in this case we need 
// an array of 1024 (1K) 32-bit elements (1024 elements where each element is 32-bit wide).  
// for example, to declare an array of 256 32-bit elements, declaration is: reg[31:0] memory[0:255]
////////////////////////////////////////////////////////////////////////////////

module DataMemory(Address, WriteData, Clk, MemWrite, MemRead, ReadData); 

    input [31:0] Address; 	// Input Address 
    input [31:0] WriteData; // Data that needs to be written into the address 
    input Clk;
    input MemWrite; 		// Control signal for memory write 
    input MemRead; 			// Control signal for memory read 

    output reg[31:0] ReadData; // Contents of memory location at Address

    // reg [31:0] memory [0:1023]; // Modified for task3
    reg [31:0] memory [0:16383];

    // Initialize Data Memory - Task2
    initial begin
	 memory[0] = 32'd4;          
     memory[1] = 32'd45;
     memory[2] = 32'd54;
     memory[3] = 32'd69;
     memory[4] = 32'd19;
     memory[5] = 32'd42;
     memory[6] = 32'd35;
     memory[7] = 32'd91;
     memory[8] = 32'd48;
     memory[9] = 32'd37;
     memory[10] = 32'd66;
     memory[11] = 32'd25;
     memory[12] = 32'd32;
     memory[13] = 32'd90;
     memory[14] = 32'd18;
     memory[15] = 32'd12;
     memory[16] = 32'd26;
     memory[17] = 32'd18;
     memory[18] = 32'd234;
     memory[19] = 32'd84;
     memory[20] = 32'd93;
     memory[21] = 32'd215;
     memory[22] = 32'd123;
     memory[23] = 32'd47;
     memory[24] = 32'd220;
     memory[25] = 32'd217;
     memory[26] = 32'd181;
     memory[27] = 32'd222;
     memory[28] = 32'd12;
     memory[29] = 32'd83;
     memory[30] = 32'd204;
     memory[31] = 32'd12;
     memory[32] = 32'd219;
     memory[33] = 32'd32;
     memory[34] = 32'd139;
     memory[35] = 32'd86;
     memory[36] = 32'd9;
     memory[37] = 32'd248;
     memory[38] = 32'd77;
     memory[39] = 32'd49;
     memory[40] = 32'd45;
     memory[41] = 32'd97;
     memory[42] = 32'd58;
     memory[43] = 32'd215;
     memory[44] = 32'd67;
     memory[45] = 32'd71;
     memory[46] = 32'd60;
     memory[47] = 32'd129;
     memory[48] = 32'd162;
     memory[49] = 32'd122;
     memory[50] = 32'd78;
     memory[51] = 32'd104;
     memory[52] = 32'd93;
     memory[53] = 32'd92;
     memory[54] = 32'd254;
     memory[55] = 32'd181;
     memory[56] = 32'd17;
     memory[57] = 32'd231;
     memory[58] = 32'd220;
     memory[59] = 32'd97;
     memory[60] = 32'd196;
     memory[61] = 32'd131;
     memory[62] = 32'd119;
     memory[63] = 32'd29;
     memory[64] = 32'd149;
     memory[65] = 32'd98;
     memory[66] = 32'd133;
     memory[67] = 32'd148;
     memory[68] = 32'd123;
     memory[69] = 32'd174;
     memory[70] = 32'd180;
     memory[71] = 32'd2;
     memory[72] = 32'd37;
     memory[73] = 32'd170;
     memory[74] = 32'd11;
     memory[75] = 32'd196;
     memory[76] = 32'd182;
     memory[77] = 32'd220;
     memory[78] = 32'd218;
     memory[79] = 32'd202;
     memory[80] = 32'd36;
     memory[81] = 32'd193;
     memory[82] = 32'd108;
     memory[83] = 32'd217;
     memory[84] = 32'd220;
     memory[85] = 32'd233;
     memory[86] = 32'd221;
     memory[87] = 32'd175;
     memory[88] = 32'd154;
     memory[89] = 32'd213;
     memory[90] = 32'd223;
     memory[91] = 32'd22;
     memory[92] = 32'd211;
     memory[93] = 32'd222;
     memory[94] = 32'd103;
     memory[95] = 32'd131;
     memory[96] = 32'd249;
     memory[97] = 32'd40;
     memory[98] = 32'd113;
     memory[99] = 32'd117;
     memory[100] = 32'd2;
     memory[101] = 32'd2;
     memory[102] = 32'd159;
     memory[103] = 32'd90;
     memory[104] = 32'd53;
     memory[105] = 32'd129;
     memory[106] = 32'd252;
     memory[107] = 32'd166;
     memory[108] = 32'd122;
     memory[109] = 32'd85;
     memory[110] = 32'd217;
     memory[111] = 32'd200;
     memory[112] = 32'd50;
     memory[113] = 32'd83;
     memory[114] = 32'd189;
     memory[115] = 32'd74;
     memory[116] = 32'd69;
     memory[117] = 32'd180;
     memory[118] = 32'd46;
     memory[119] = 32'd2;
     memory[120] = 32'd216;
     memory[121] = 32'd123;
     memory[122] = 32'd244;
     memory[123] = 32'd253;
     memory[124] = 32'd229;
     memory[125] = 32'd63;
     memory[126] = 32'd48;
     memory[127] = 32'd219;
     memory[128] = 32'd66;
     memory[129] = 32'd218;
     memory[130] = 32'd40;
     memory[131] = 32'd25;
     memory[132] = 32'd212;
     memory[133] = 32'd12;
     memory[134] = 32'd194;
     memory[135] = 32'd152;
     memory[136] = 32'd130;
     memory[137] = 32'd181;
     memory[138] = 32'd215;
     memory[139] = 32'd158;
     memory[140] = 32'd132;
     memory[141] = 32'd124;
     memory[142] = 32'd100;
     memory[143] = 32'd28;
     memory[144] = 32'd190;
     memory[145] = 32'd41;
     memory[146] = 32'd35;
     memory[147] = 32'd141;
     memory[148] = 32'd4;
     memory[149] = 32'd69;
     memory[150] = 32'd89;
     memory[151] = 32'd16;
     memory[152] = 32'd230;
     memory[153] = 32'd23;
     memory[154] = 32'd43;
     memory[155] = 32'd245;
     memory[156] = 32'd148;
     memory[157] = 32'd80;
     memory[158] = 32'd150;
     memory[159] = 32'd99;
     memory[160] = 32'd126;
     memory[161] = 32'd114;
     memory[162] = 32'd215;
     memory[163] = 32'd53;
     memory[164] = 32'd205;
     memory[165] = 32'd114;
     memory[166] = 32'd162;
     memory[167] = 32'd231;
     memory[168] = 32'd75;
     memory[169] = 32'd66;
     memory[170] = 32'd102;
     memory[171] = 32'd192;
     memory[172] = 32'd134;
     memory[173] = 32'd173;
     memory[174] = 32'd128;
     memory[175] = 32'd202;
     memory[176] = 32'd106;
     memory[177] = 32'd148;
     memory[178] = 32'd132;
     memory[179] = 32'd103;
     memory[180] = 32'd164;
     memory[181] = 32'd224;
     memory[182] = 32'd101;
     memory[183] = 32'd8;
     memory[184] = 32'd7;
     memory[185] = 32'd24;
     memory[186] = 32'd13;
     memory[187] = 32'd41;
     memory[188] = 32'd19;
     memory[189] = 32'd166;
     memory[190] = 32'd46;
     memory[191] = 32'd188;
     memory[192] = 32'd226;
     memory[193] = 32'd78;
     memory[194] = 32'd192;
     memory[195] = 32'd42;
     memory[196] = 32'd17;
     memory[197] = 32'd146;
     memory[198] = 32'd243;
     memory[199] = 32'd171;
     memory[200] = 32'd46;
     memory[201] = 32'd14;
     memory[202] = 32'd81;
     memory[203] = 32'd68;
     memory[204] = 32'd159;
     memory[205] = 32'd129;
     memory[206] = 32'd251;
     memory[207] = 32'd27;
     memory[208] = 32'd99;
     memory[209] = 32'd130;
     memory[210] = 32'd185;
     memory[211] = 32'd143;
     memory[212] = 32'd95;
     memory[213] = 32'd20;
     memory[214] = 32'd93;
     memory[215] = 32'd236;
     memory[216] = 32'd154;
     memory[217] = 32'd234;
     memory[218] = 32'd155;
     memory[219] = 32'd246;
     memory[220] = 32'd187;
     memory[221] = 32'd117;
     memory[222] = 32'd189;
     memory[223] = 32'd89;
     memory[224] = 32'd135;
     memory[225] = 32'd194;
     memory[226] = 32'd108;
     memory[227] = 32'd104;
     memory[228] = 32'd50;
     memory[229] = 32'd168;
     memory[230] = 32'd90;
     memory[231] = 32'd35;
     memory[232] = 32'd119;
     memory[233] = 32'd184;
     memory[234] = 32'd207;
     memory[235] = 32'd232;
     memory[236] = 32'd238;
     memory[237] = 32'd22;
     memory[238] = 32'd188;
     memory[239] = 32'd18;
     memory[240] = 32'd25;
     memory[241] = 32'd203;
     memory[242] = 32'd157;
     memory[243] = 32'd180;
     memory[244] = 32'd168;
     memory[245] = 32'd2;
     memory[246] = 32'd202;
     memory[247] = 32'd238;
     memory[248] = 32'd118;
     memory[249] = 32'd176;
     memory[250] = 32'd203;
     memory[251] = 32'd207;
     memory[252] = 32'd96;
     memory[253] = 32'd247;
     memory[254] = 32'd218;
     memory[255] = 32'd100;
     memory[256] = 32'd150;
     memory[257] = 32'd151;
     memory[258] = 32'd252;
     memory[259] = 32'd75;
     memory[260] = 32'd147;
     memory[261] = 32'd79;
     memory[262] = 32'd217;
     memory[263] = 32'd19;
     memory[264] = 32'd160;
     memory[265] = 32'd194;
     memory[266] = 32'd89;
     memory[267] = 32'd162;
     memory[268] = 32'd18;
     memory[269] = 32'd241;
     memory[270] = 32'd10;
     memory[271] = 32'd80;
     memory[272] = 32'd103;
     memory[273] = 32'd75;
     memory[274] = 32'd180;
     memory[275] = 32'd34;
     memory[276] = 32'd149;
     memory[277] = 32'd75;
     memory[278] = 32'd47;
     memory[279] = 32'd223;
     memory[280] = 32'd30;
     memory[281] = 32'd6;
     memory[282] = 32'd32;
     memory[283] = 32'd210;
     memory[284] = 32'd187;
     memory[285] = 32'd179;
     memory[286] = 32'd16;
     memory[287] = 32'd225;
     memory[288] = 32'd101;
     memory[289] = 32'd150;
     memory[290] = 32'd233;
     memory[291] = 32'd254;
     memory[292] = 32'd236;
     memory[293] = 32'd78;
     memory[294] = 32'd238;
     memory[295] = 32'd167;
     memory[296] = 32'd21;
     memory[297] = 32'd195;
     memory[298] = 32'd172;
     memory[299] = 32'd18;
     memory[300] = 32'd57;
     memory[301] = 32'd151;
     memory[302] = 32'd24;
     memory[303] = 32'd20;
     memory[304] = 32'd55;
     memory[305] = 32'd200;
     memory[306] = 32'd46;
     memory[307] = 32'd61;
     memory[308] = 32'd108;
     memory[309] = 32'd149;
     memory[310] = 32'd186;
     memory[311] = 32'd17;
     memory[312] = 32'd10;
     memory[313] = 32'd110;
     memory[314] = 32'd226;
     memory[315] = 32'd118;
     memory[316] = 32'd128;
     memory[317] = 32'd109;
     memory[318] = 32'd27;
     memory[319] = 32'd152;
     memory[320] = 32'd124;
     memory[321] = 32'd217;
     memory[322] = 32'd123;
     memory[323] = 32'd210;
     memory[324] = 32'd112;
     memory[325] = 32'd92;
     memory[326] = 32'd130;
     memory[327] = 32'd174;
     memory[328] = 32'd4;
     memory[329] = 32'd95;
     memory[330] = 32'd28;
     memory[331] = 32'd85;
     memory[332] = 32'd130;
     memory[333] = 32'd175;
     memory[334] = 32'd53;
     memory[335] = 32'd121;
     memory[336] = 32'd72;
     memory[337] = 32'd45;
     memory[338] = 32'd68;
     memory[339] = 32'd105;
     memory[340] = 32'd183;
     memory[341] = 32'd193;
     memory[342] = 32'd23;
     memory[343] = 32'd120;
     memory[344] = 32'd23;
     memory[345] = 32'd204;
     memory[346] = 32'd169;
     memory[347] = 32'd51;
     memory[348] = 32'd37;
     memory[349] = 32'd71;
     memory[350] = 32'd178;
     memory[351] = 32'd69;
     memory[352] = 32'd186;
     memory[353] = 32'd140;
     memory[354] = 32'd198;
     memory[355] = 32'd198;
     memory[356] = 32'd7;
     memory[357] = 32'd174;
     memory[358] = 32'd175;
     memory[359] = 32'd143;
     memory[360] = 32'd223;
     memory[361] = 32'd67;
     memory[362] = 32'd184;
     memory[363] = 32'd245;
     memory[364] = 32'd229;
     memory[365] = 32'd22;
     memory[366] = 32'd74;
     memory[367] = 32'd14;
     memory[368] = 32'd162;
     memory[369] = 32'd40;
     memory[370] = 32'd56;
     memory[371] = 32'd69;
     memory[372] = 32'd78;
     memory[373] = 32'd43;
     memory[374] = 32'd48;
     memory[375] = 32'd11;
     memory[376] = 32'd246;
     memory[377] = 32'd121;
     memory[378] = 32'd19;
     memory[379] = 32'd124;
     memory[380] = 32'd221;
     memory[381] = 32'd72;
     memory[382] = 32'd86;
     memory[383] = 32'd201;
     memory[384] = 32'd138;
     memory[385] = 32'd91;
     memory[386] = 32'd110;
     memory[387] = 32'd5;
     memory[388] = 32'd159;
     memory[389] = 32'd29;
     memory[390] = 32'd89;
     memory[391] = 32'd12;
     memory[392] = 32'd162;
     memory[393] = 32'd116;
     memory[394] = 32'd56;
     memory[395] = 32'd101;
     memory[396] = 32'd145;
     memory[397] = 32'd218;
     memory[398] = 32'd114;
     memory[399] = 32'd221;
     memory[400] = 32'd57;
     memory[401] = 32'd8;
     memory[402] = 32'd205;
     memory[403] = 32'd80;
     memory[404] = 32'd147;
     memory[405] = 32'd165;
     memory[406] = 32'd164;
     memory[407] = 32'd240;
     memory[408] = 32'd196;
     memory[409] = 32'd23;
     memory[410] = 32'd235;
     memory[411] = 32'd97;
     memory[412] = 32'd233;
     memory[413] = 32'd105;
     memory[414] = 32'd165;
     memory[415] = 32'd185;
     memory[416] = 32'd43;
     memory[417] = 32'd79;
     memory[418] = 32'd197;
     memory[419] = 32'd4;
     memory[420] = 32'd126;
     memory[421] = 32'd221;
     memory[422] = 32'd226;
     memory[423] = 32'd52;
     memory[424] = 32'd65;
     memory[425] = 32'd8;
     memory[426] = 32'd127;
     memory[427] = 32'd163;
     memory[428] = 32'd9;
     memory[429] = 32'd29;
     memory[430] = 32'd176;
     memory[431] = 32'd219;
     memory[432] = 32'd96;
     memory[433] = 32'd201;
     memory[434] = 32'd126;
     memory[435] = 32'd146;
     memory[436] = 32'd211;
     memory[437] = 32'd77;
     memory[438] = 32'd159;
     memory[439] = 32'd200;
     memory[440] = 32'd81;
     memory[441] = 32'd147;
     memory[442] = 32'd111;
     memory[443] = 32'd253;
     memory[444] = 32'd224;
     memory[445] = 32'd6;
     memory[446] = 32'd228;
     memory[447] = 32'd205;
     memory[448] = 32'd115;
     memory[449] = 32'd29;
     memory[450] = 32'd221;
     memory[451] = 32'd220;
     memory[452] = 32'd172;
     memory[453] = 32'd25;
     memory[454] = 32'd188;
     memory[455] = 32'd109;
     memory[456] = 32'd117;
     memory[457] = 32'd210;
     memory[458] = 32'd113;
     memory[459] = 32'd220;
     memory[460] = 32'd241;
     memory[461] = 32'd248;
     memory[462] = 32'd46;
     memory[463] = 32'd4;
     memory[464] = 32'd23;
     memory[465] = 32'd62;
     memory[466] = 32'd201;
     memory[467] = 32'd184;
     memory[468] = 32'd167;
     memory[469] = 32'd90;
     memory[470] = 32'd72;
     memory[471] = 32'd194;
     memory[472] = 32'd130;
     memory[473] = 32'd223;
     memory[474] = 32'd45;
     memory[475] = 32'd98;
     memory[476] = 32'd227;
     memory[477] = 32'd27;
     memory[478] = 32'd11;
     memory[479] = 32'd8;
     memory[480] = 32'd211;
     memory[481] = 32'd163;
     memory[482] = 32'd126;
     memory[483] = 32'd116;
     memory[484] = 32'd230;
     memory[485] = 32'd63;
     memory[486] = 32'd1;
     memory[487] = 32'd177;
     memory[488] = 32'd155;
     memory[489] = 32'd69;
     memory[490] = 32'd174;
     memory[491] = 32'd143;
     memory[492] = 32'd101;
     memory[493] = 32'd3;
     memory[494] = 32'd143;
     memory[495] = 32'd212;
     memory[496] = 32'd67;
     memory[497] = 32'd79;
     memory[498] = 32'd99;
     memory[499] = 32'd10;
     memory[500] = 32'd104;
     memory[501] = 32'd140;
     memory[502] = 32'd57;
     memory[503] = 32'd186;
     memory[504] = 32'd214;
     memory[505] = 32'd69;
     memory[506] = 32'd174;
     memory[507] = 32'd199;
     memory[508] = 32'd71;
     memory[509] = 32'd98;
     memory[510] = 32'd172;
     memory[511] = 32'd146;
     memory[512] = 32'd5;
     memory[513] = 32'd221;
     memory[514] = 32'd89;
     memory[515] = 32'd245;
     memory[516] = 32'd209;
     memory[517] = 32'd80;
     memory[518] = 32'd147;
     memory[519] = 32'd100;
     memory[520] = 32'd230;
     memory[521] = 32'd108;
     memory[522] = 32'd111;
     memory[523] = 32'd95;
     memory[524] = 32'd249;
     memory[525] = 32'd214;
     memory[526] = 32'd4;
     memory[527] = 32'd56;
     memory[528] = 32'd84;
     memory[529] = 32'd43;
     memory[530] = 32'd162;
     memory[531] = 32'd104;
     memory[532] = 32'd149;
     memory[533] = 32'd77;
     memory[534] = 32'd238;
     memory[535] = 32'd28;
     memory[536] = 32'd165;
     memory[537] = 32'd9;
     memory[538] = 32'd220;
     memory[539] = 32'd172;
     memory[540] = 32'd225;
     memory[541] = 32'd210;
     memory[542] = 32'd21;
     memory[543] = 32'd219;
     memory[544] = 32'd175;
     memory[545] = 32'd233;
     memory[546] = 32'd170;
     memory[547] = 32'd92;
     memory[548] = 32'd133;
     memory[549] = 32'd23;
     memory[550] = 32'd58;
     memory[551] = 32'd109;
     memory[552] = 32'd243;
     memory[553] = 32'd137;
     memory[554] = 32'd240;
     memory[555] = 32'd157;
     memory[556] = 32'd64;
     memory[557] = 32'd216;
     memory[558] = 32'd14;
     memory[559] = 32'd4;
     memory[560] = 32'd71;
     memory[561] = 32'd176;
     memory[562] = 32'd165;
     memory[563] = 32'd90;
     memory[564] = 32'd104;
     memory[565] = 32'd65;
     memory[566] = 32'd143;
     memory[567] = 32'd180;
     memory[568] = 32'd63;
     memory[569] = 32'd37;
     memory[570] = 32'd43;
     memory[571] = 32'd0;
     memory[572] = 32'd5;
     memory[573] = 32'd211;
     memory[574] = 32'd189;
     memory[575] = 32'd143;
     memory[576] = 32'd91;
     memory[577] = 32'd223;
     memory[578] = 32'd219;
     memory[579] = 32'd216;
     memory[580] = 32'd21;
     memory[581] = 32'd202;
     memory[582] = 32'd76;
     memory[583] = 32'd107;
     memory[584] = 32'd69;
     memory[585] = 32'd190;
     memory[586] = 32'd176;
     memory[587] = 32'd109;
     memory[588] = 32'd42;
     memory[589] = 32'd143;
     memory[590] = 32'd250;
     memory[591] = 32'd116;
     memory[592] = 32'd35;
     memory[593] = 32'd12;
     memory[594] = 32'd214;
     memory[595] = 32'd190;
     memory[596] = 32'd189;
     memory[597] = 32'd172;
     memory[598] = 32'd141;
     memory[599] = 32'd105;
     memory[600] = 32'd80;
     memory[601] = 32'd112;
     memory[602] = 32'd118;
     memory[603] = 32'd52;
     memory[604] = 32'd10;
     memory[605] = 32'd65;
     memory[606] = 32'd44;
     memory[607] = 32'd236;
     memory[608] = 32'd235;
     memory[609] = 32'd18;
     memory[610] = 32'd157;
     memory[611] = 32'd159;
     memory[612] = 32'd184;
     memory[613] = 32'd122;
     memory[614] = 32'd214;
     memory[615] = 32'd251;
     memory[616] = 32'd244;
     memory[617] = 32'd57;
     memory[618] = 32'd20;
     memory[619] = 32'd238;
     memory[620] = 32'd71;
     memory[621] = 32'd28;
     memory[622] = 32'd36;
     memory[623] = 32'd231;
     memory[624] = 32'd101;
     memory[625] = 32'd53;
     memory[626] = 32'd189;
     memory[627] = 32'd72;
     memory[628] = 32'd126;
     memory[629] = 32'd11;
     memory[630] = 32'd78;
     memory[631] = 32'd208;
     memory[632] = 32'd17;
     memory[633] = 32'd172;
     memory[634] = 32'd133;
     memory[635] = 32'd202;
     memory[636] = 32'd95;
     memory[637] = 32'd32;
     memory[638] = 32'd200;
     memory[639] = 32'd44;
     memory[640] = 32'd93;
     memory[641] = 32'd230;
     memory[642] = 32'd62;
     memory[643] = 32'd29;
     memory[644] = 32'd23;
     memory[645] = 32'd92;
     memory[646] = 32'd114;
     memory[647] = 32'd205;
     memory[648] = 32'd226;
     memory[649] = 32'd251;
     memory[650] = 32'd29;
     memory[651] = 32'd167;
     memory[652] = 32'd172;
     memory[653] = 32'd15;
     memory[654] = 32'd92;
     memory[655] = 32'd36;
     memory[656] = 32'd250;
     memory[657] = 32'd197;
     memory[658] = 32'd175;
     memory[659] = 32'd235;
     memory[660] = 32'd64;
     memory[661] = 32'd204;
     memory[662] = 32'd213;
     memory[663] = 32'd136;
     memory[664] = 32'd148;
     memory[665] = 32'd110;
     memory[666] = 32'd131;
     memory[667] = 32'd154;
     memory[668] = 32'd91;
     memory[669] = 32'd108;
     memory[670] = 32'd131;
     memory[671] = 32'd186;
     memory[672] = 32'd156;
     memory[673] = 32'd54;
     memory[674] = 32'd202;
     memory[675] = 32'd49;
     memory[676] = 32'd121;
     memory[677] = 32'd75;
     memory[678] = 32'd161;
     memory[679] = 32'd244;
     memory[680] = 32'd201;
     memory[681] = 32'd218;
     memory[682] = 32'd171;
     memory[683] = 32'd239;
     memory[684] = 32'd183;
     memory[685] = 32'd114;
     memory[686] = 32'd41;
     memory[687] = 32'd126;
     memory[688] = 32'd229;
     memory[689] = 32'd15;
     memory[690] = 32'd56;
     memory[691] = 32'd5;
     memory[692] = 32'd248;
     memory[693] = 32'd220;
     memory[694] = 32'd41;
     memory[695] = 32'd146;
     memory[696] = 32'd155;
     memory[697] = 32'd137;
     memory[698] = 32'd141;
     memory[699] = 32'd213;
     memory[700] = 32'd253;
     memory[701] = 32'd72;
     memory[702] = 32'd240;
     memory[703] = 32'd59;
     memory[704] = 32'd55;
     memory[705] = 32'd248;
     memory[706] = 32'd71;
     memory[707] = 32'd198;
     memory[708] = 32'd71;
     memory[709] = 32'd134;
     memory[710] = 32'd24;
     memory[711] = 32'd221;
     memory[712] = 32'd38;
     memory[713] = 32'd83;
     memory[714] = 32'd33;
     memory[715] = 32'd136;
     memory[716] = 32'd4;
     memory[717] = 32'd121;
     memory[718] = 32'd134;
     memory[719] = 32'd42;
     memory[720] = 32'd106;
     memory[721] = 32'd168;
     memory[722] = 32'd105;
     memory[723] = 32'd205;
     memory[724] = 32'd46;
     memory[725] = 32'd228;
     memory[726] = 32'd97;
     memory[727] = 32'd35;
     memory[728] = 32'd56;
     memory[729] = 32'd173;
     memory[730] = 32'd8;
     memory[731] = 32'd76;
     memory[732] = 32'd159;
     memory[733] = 32'd132;
     memory[734] = 32'd207;
     memory[735] = 32'd13;
     memory[736] = 32'd26;
     memory[737] = 32'd206;
     memory[738] = 32'd23;
     memory[739] = 32'd235;
     memory[740] = 32'd43;
     memory[741] = 32'd249;
     memory[742] = 32'd121;
     memory[743] = 32'd104;
     memory[744] = 32'd20;
     memory[745] = 32'd109;
     memory[746] = 32'd19;
     memory[747] = 32'd35;
     memory[748] = 32'd172;
     memory[749] = 32'd165;
     memory[750] = 32'd25;
     memory[751] = 32'd147;
     memory[752] = 32'd196;
     memory[753] = 32'd126;
     memory[754] = 32'd36;
     memory[755] = 32'd191;
     memory[756] = 32'd162;
     memory[757] = 32'd29;
     memory[758] = 32'd66;
     memory[759] = 32'd117;
     memory[760] = 32'd233;
     memory[761] = 32'd130;
     memory[762] = 32'd252;
     memory[763] = 32'd132;
     memory[764] = 32'd244;
     memory[765] = 32'd170;
     memory[766] = 32'd153;
     memory[767] = 32'd46;
     memory[768] = 32'd205;
     memory[769] = 32'd9;
     memory[770] = 32'd156;
     memory[771] = 32'd163;
     memory[772] = 32'd201;
     memory[773] = 32'd5;
     memory[774] = 32'd78;
     memory[775] = 32'd214;
     memory[776] = 32'd26;
     memory[777] = 32'd195;
     memory[778] = 32'd187;
     memory[779] = 32'd82;
     memory[780] = 32'd105;
     memory[781] = 32'd101;
     memory[782] = 32'd230;
     memory[783] = 32'd25;
     memory[784] = 32'd150;
     memory[785] = 32'd32;
     memory[786] = 32'd57;
     memory[787] = 32'd118;
     memory[788] = 32'd221;
     memory[789] = 32'd144;
     memory[790] = 32'd53;
     memory[791] = 32'd181;
     memory[792] = 32'd35;
     memory[793] = 32'd242;
     memory[794] = 32'd111;
     memory[795] = 32'd101;
     memory[796] = 32'd150;
     memory[797] = 32'd36;
     memory[798] = 32'd246;
     memory[799] = 32'd236;
     memory[800] = 32'd98;
     memory[801] = 32'd14;
     memory[802] = 32'd69;
     memory[803] = 32'd64;
     memory[804] = 32'd86;
     memory[805] = 32'd1;
     memory[806] = 32'd159;
     memory[807] = 32'd185;
     memory[808] = 32'd210;
     memory[809] = 32'd191;
     memory[810] = 32'd222;
     memory[811] = 32'd34;
     memory[812] = 32'd161;
     memory[813] = 32'd5;
     memory[814] = 32'd100;
     memory[815] = 32'd192;
     memory[816] = 32'd98;
     memory[817] = 32'd54;
     memory[818] = 32'd7;
     memory[819] = 32'd165;
     memory[820] = 32'd17;
     memory[821] = 32'd248;
     memory[822] = 32'd235;
     memory[823] = 32'd30;
     memory[824] = 32'd98;
     memory[825] = 32'd73;
     memory[826] = 32'd41;
     memory[827] = 32'd150;
     memory[828] = 32'd13;
     memory[829] = 32'd40;
     memory[830] = 32'd192;
     memory[831] = 32'd101;
     memory[832] = 32'd75;
     memory[833] = 32'd153;
     memory[834] = 32'd191;
     memory[835] = 32'd175;
     memory[836] = 32'd121;
     memory[837] = 32'd217;
     memory[838] = 32'd180;
     memory[839] = 32'd2;
     memory[840] = 32'd25;
     memory[841] = 32'd61;
     memory[842] = 32'd104;
     memory[843] = 32'd57;
     memory[844] = 32'd175;
     memory[845] = 32'd19;
     memory[846] = 32'd89;
     memory[847] = 32'd193;
     memory[848] = 32'd134;
     memory[849] = 32'd207;
     memory[850] = 32'd10;
     memory[851] = 32'd28;
     memory[852] = 32'd83;
     memory[853] = 32'd226;
     memory[854] = 32'd201;
     memory[855] = 32'd50;
     memory[856] = 32'd125;
     memory[857] = 32'd135;
     memory[858] = 32'd152;
     memory[859] = 32'd111;
     memory[860] = 32'd44;
     memory[861] = 32'd144;
     memory[862] = 32'd98;
     memory[863] = 32'd183;
     memory[864] = 32'd195;
     memory[865] = 32'd215;
     memory[866] = 32'd19;
     memory[867] = 32'd39;
     memory[868] = 32'd52;
     memory[869] = 32'd173;
     memory[870] = 32'd0;
     memory[871] = 32'd106;
     memory[872] = 32'd229;
     memory[873] = 32'd238;
     memory[874] = 32'd137;
     memory[875] = 32'd205;
     memory[876] = 32'd84;
     memory[877] = 32'd99;
     memory[878] = 32'd213;
     memory[879] = 32'd122;
     memory[880] = 32'd72;
     memory[881] = 32'd95;
     memory[882] = 32'd94;
     memory[883] = 32'd12;
     memory[884] = 32'd134;
     memory[885] = 32'd180;
     memory[886] = 32'd207;
     memory[887] = 32'd194;
     memory[888] = 32'd166;
     memory[889] = 32'd57;
     memory[890] = 32'd17;
     memory[891] = 32'd87;
     memory[892] = 32'd42;
     memory[893] = 32'd164;
     memory[894] = 32'd158;
     memory[895] = 32'd184;
     memory[896] = 32'd109;
     memory[897] = 32'd187;
     memory[898] = 32'd152;
     memory[899] = 32'd226;
     memory[900] = 32'd57;
     memory[901] = 32'd94;
     memory[902] = 32'd136;
     memory[903] = 32'd209;
     memory[904] = 32'd86;
     memory[905] = 32'd3;
     memory[906] = 32'd79;
     memory[907] = 32'd71;
     memory[908] = 32'd175;
     memory[909] = 32'd72;
     memory[910] = 32'd71;
     memory[911] = 32'd34;
     memory[912] = 32'd59;
     memory[913] = 32'd72;
     memory[914] = 32'd48;
     memory[915] = 32'd247;
     memory[916] = 32'd174;
     memory[917] = 32'd77;
     memory[918] = 32'd157;
     memory[919] = 32'd220;
     memory[920] = 32'd133;
     memory[921] = 32'd22;
     memory[922] = 32'd109;
     memory[923] = 32'd212;
     memory[924] = 32'd56;
     memory[925] = 32'd254;
     memory[926] = 32'd217;
     memory[927] = 32'd37;
     memory[928] = 32'd236;
     memory[929] = 32'd74;
     memory[930] = 32'd184;
     memory[931] = 32'd75;
     memory[932] = 32'd79;
     memory[933] = 32'd171;
     memory[934] = 32'd37;
     memory[935] = 32'd62;
     memory[936] = 32'd44;
     memory[937] = 32'd24;
     memory[938] = 32'd149;
     memory[939] = 32'd26;
     memory[940] = 32'd201;
     memory[941] = 32'd90;
     memory[942] = 32'd2;
     memory[943] = 32'd166;
     memory[944] = 32'd236;
     memory[945] = 32'd63;
     memory[946] = 32'd64;
     memory[947] = 32'd73;
     memory[948] = 32'd106;
     memory[949] = 32'd52;
     memory[950] = 32'd45;
     memory[951] = 32'd33;
     memory[952] = 32'd82;
     memory[953] = 32'd88;
     memory[954] = 32'd105;
     memory[955] = 32'd131;
     memory[956] = 32'd95;
     memory[957] = 32'd40;
     memory[958] = 32'd32;
     memory[959] = 32'd39;
     memory[960] = 32'd214;
     memory[961] = 32'd179;
     memory[962] = 32'd69;
     memory[963] = 32'd52;
     memory[964] = 32'd233;
     memory[965] = 32'd109;
     memory[966] = 32'd228;
     memory[967] = 32'd39;
     memory[968] = 32'd9;
     memory[969] = 32'd104;
     memory[970] = 32'd18;
     memory[971] = 32'd54;
     memory[972] = 32'd165;
     memory[973] = 32'd164;
     memory[974] = 32'd155;
     memory[975] = 32'd96;
     memory[976] = 32'd43;
     memory[977] = 32'd234;
     memory[978] = 32'd50;
     memory[979] = 32'd106;
     memory[980] = 32'd124;
     memory[981] = 32'd2;
     memory[982] = 32'd21;
     memory[983] = 32'd164;
     memory[984] = 32'd167;
     memory[985] = 32'd168;
     memory[986] = 32'd40;
     memory[987] = 32'd251;
     memory[988] = 32'd147;
     memory[989] = 32'd15;
     memory[990] = 32'd201;
     memory[991] = 32'd137;
     memory[992] = 32'd59;
     memory[993] = 32'd29;
     memory[994] = 32'd124;
     memory[995] = 32'd50;
     memory[996] = 32'd207;
     memory[997] = 32'd36;
     memory[998] = 32'd134;
     memory[999] = 32'd107;
     memory[1000] = 32'd107;
     memory[1001] = 32'd160;
     memory[1002] = 32'd52;
     memory[1003] = 32'd220;
     memory[1004] = 32'd253;
     memory[1005] = 32'd86;
     memory[1006] = 32'd234;
     memory[1007] = 32'd245;
     memory[1008] = 32'd6;
     memory[1009] = 32'd103;
     memory[1010] = 32'd56;
     memory[1011] = 32'd168;
     memory[1012] = 32'd152;
     memory[1013] = 32'd189;
     memory[1014] = 32'd42;
     memory[1015] = 32'd215;
     memory[1016] = 32'd81;
     memory[1017] = 32'd54;
     memory[1018] = 32'd130;
     memory[1019] = 32'd138;
     memory[1020] = 32'd60;
     memory[1021] = 32'd235;
     memory[1022] = 32'd141;
     memory[1023] = 32'd227;
     memory[1024] = 32'd134;
     memory[1025] = 32'd124;
     memory[1026] = 32'd0;
     memory[1027] = 32'd224;
     memory[1028] = 32'd131;
     memory[1029] = 32'd127;
     memory[1030] = 32'd100;
     memory[1031] = 32'd249;
     memory[1032] = 32'd244;
     memory[1033] = 32'd140;
     memory[1034] = 32'd30;
     memory[1035] = 32'd144;
     memory[1036] = 32'd215;
     memory[1037] = 32'd42;
     memory[1038] = 32'd58;
     memory[1039] = 32'd237;
     memory[1040] = 32'd193;
     memory[1041] = 32'd172;
     memory[1042] = 32'd169;
     memory[1043] = 32'd221;
     memory[1044] = 32'd205;
     memory[1045] = 32'd238;
     memory[1046] = 32'd143;
     memory[1047] = 32'd247;
     memory[1048] = 32'd61;
     memory[1049] = 32'd244;
     memory[1050] = 32'd144;
     memory[1051] = 32'd74;
     memory[1052] = 32'd139;
     memory[1053] = 32'd15;
     memory[1054] = 32'd128;
     memory[1055] = 32'd102;
     memory[1056] = 32'd244;
     memory[1057] = 32'd84;
     memory[1058] = 32'd12;
     memory[1059] = 32'd127;
     memory[1060] = 32'd28;
     memory[1061] = 32'd86;
     memory[1062] = 32'd178;
     memory[1063] = 32'd8;
     memory[1064] = 32'd184;
     memory[1065] = 32'd1;
     memory[1066] = 32'd210;
     memory[1067] = 32'd186;
     memory[1068] = 32'd224;
     memory[1069] = 32'd144;
     memory[1070] = 32'd174;
     memory[1071] = 32'd131;
     memory[1072] = 32'd171;
     memory[1073] = 32'd244;
     memory[1074] = 32'd145;
     memory[1075] = 32'd101;
     memory[1076] = 32'd97;
     memory[1077] = 32'd253;
     memory[1078] = 32'd129;
     memory[1079] = 32'd227;
     memory[1080] = 32'd56;
     memory[1081] = 32'd159;
     memory[1082] = 32'd244;
     memory[1083] = 32'd13;
     memory[1084] = 32'd138;
     memory[1085] = 32'd245;
     memory[1086] = 32'd249;
     memory[1087] = 32'd147;
     memory[1088] = 32'd88;
     memory[1089] = 32'd172;
     memory[1090] = 32'd69;
     memory[1091] = 32'd127;
     memory[1092] = 32'd17;
     memory[1093] = 32'd160;
     memory[1094] = 32'd4;
     memory[1095] = 32'd46;
     memory[1096] = 32'd92;
     memory[1097] = 32'd118;
     memory[1098] = 32'd248;
     memory[1099] = 32'd34;
     memory[1100] = 32'd172;
     memory[1101] = 32'd14;
     memory[1102] = 32'd92;
     memory[1103] = 32'd72;
     memory[1104] = 32'd125;
     memory[1105] = 32'd80;
     memory[1106] = 32'd186;
     memory[1107] = 32'd178;
     memory[1108] = 32'd235;
     memory[1109] = 32'd215;
     memory[1110] = 32'd57;
     memory[1111] = 32'd34;
     memory[1112] = 32'd30;
     memory[1113] = 32'd84;
     memory[1114] = 32'd219;
     memory[1115] = 32'd116;
     memory[1116] = 32'd222;
     memory[1117] = 32'd18;
     memory[1118] = 32'd149;
     memory[1119] = 32'd45;
     memory[1120] = 32'd75;
     memory[1121] = 32'd92;
     memory[1122] = 32'd104;
     memory[1123] = 32'd132;
     memory[1124] = 32'd68;
     memory[1125] = 32'd120;
     memory[1126] = 32'd86;
     memory[1127] = 32'd188;
     memory[1128] = 32'd153;
     memory[1129] = 32'd168;
     memory[1130] = 32'd54;
     memory[1131] = 32'd4;
     memory[1132] = 32'd254;
     memory[1133] = 32'd212;
     memory[1134] = 32'd173;
     memory[1135] = 32'd195;
     memory[1136] = 32'd131;
     memory[1137] = 32'd89;
     memory[1138] = 32'd140;
     memory[1139] = 32'd109;
     memory[1140] = 32'd111;
     memory[1141] = 32'd136;
     memory[1142] = 32'd106;
     memory[1143] = 32'd181;
     memory[1144] = 32'd184;
     memory[1145] = 32'd115;
     memory[1146] = 32'd9;
     memory[1147] = 32'd41;
     memory[1148] = 32'd248;
     memory[1149] = 32'd247;
     memory[1150] = 32'd47;
     memory[1151] = 32'd79;
     memory[1152] = 32'd51;
     memory[1153] = 32'd173;
     memory[1154] = 32'd45;
     memory[1155] = 32'd58;
     memory[1156] = 32'd115;
     memory[1157] = 32'd153;
     memory[1158] = 32'd138;
     memory[1159] = 32'd127;
     memory[1160] = 32'd147;
     memory[1161] = 32'd20;
     memory[1162] = 32'd81;
     memory[1163] = 32'd172;
     memory[1164] = 32'd199;
     memory[1165] = 32'd244;
     memory[1166] = 32'd211;
     memory[1167] = 32'd60;
     memory[1168] = 32'd18;
     memory[1169] = 32'd3;
     memory[1170] = 32'd100;
     memory[1171] = 32'd7;
     memory[1172] = 32'd9;
     memory[1173] = 32'd90;
     memory[1174] = 32'd118;
     memory[1175] = 32'd237;
     memory[1176] = 32'd223;
     memory[1177] = 32'd154;
     memory[1178] = 32'd108;
     memory[1179] = 32'd32;
     memory[1180] = 32'd174;
     memory[1181] = 32'd111;
     memory[1182] = 32'd217;
     memory[1183] = 32'd204;
     memory[1184] = 32'd104;
     memory[1185] = 32'd245;
     memory[1186] = 32'd170;
     memory[1187] = 32'd99;
     memory[1188] = 32'd48;
     memory[1189] = 32'd223;
     memory[1190] = 32'd217;
     memory[1191] = 32'd217;
     memory[1192] = 32'd156;
     memory[1193] = 32'd83;
     memory[1194] = 32'd90;
     memory[1195] = 32'd196;
     memory[1196] = 32'd80;
     memory[1197] = 32'd61;
     memory[1198] = 32'd19;
     memory[1199] = 32'd35;
     memory[1200] = 32'd17;
     memory[1201] = 32'd69;
     memory[1202] = 32'd92;
     memory[1203] = 32'd85;
     memory[1204] = 32'd199;
     memory[1205] = 32'd49;
     memory[1206] = 32'd101;
     memory[1207] = 32'd112;
     memory[1208] = 32'd200;
     memory[1209] = 32'd29;
     memory[1210] = 32'd178;
     memory[1211] = 32'd41;
     memory[1212] = 32'd145;
     memory[1213] = 32'd88;
     memory[1214] = 32'd223;
     memory[1215] = 32'd91;
     memory[1216] = 32'd163;
     memory[1217] = 32'd126;
     memory[1218] = 32'd113;
     memory[1219] = 32'd110;
     memory[1220] = 32'd166;
     memory[1221] = 32'd213;
     memory[1222] = 32'd72;
     memory[1223] = 32'd128;
     memory[1224] = 32'd118;
     memory[1225] = 32'd7;
     memory[1226] = 32'd100;
     memory[1227] = 32'd220;
     memory[1228] = 32'd109;
     memory[1229] = 32'd125;
     memory[1230] = 32'd29;
     memory[1231] = 32'd62;
     memory[1232] = 32'd195;
     memory[1233] = 32'd197;
     memory[1234] = 32'd129;
     memory[1235] = 32'd209;
     memory[1236] = 32'd14;
     memory[1237] = 32'd95;
     memory[1238] = 32'd45;
     memory[1239] = 32'd246;
     memory[1240] = 32'd15;
     memory[1241] = 32'd115;
     memory[1242] = 32'd87;
     memory[1243] = 32'd38;
     memory[1244] = 32'd232;
     memory[1245] = 32'd184;
     memory[1246] = 32'd14;
     memory[1247] = 32'd97;
     memory[1248] = 32'd67;
     memory[1249] = 32'd13;
     memory[1250] = 32'd101;
     memory[1251] = 32'd21;
     memory[1252] = 32'd61;
     memory[1253] = 32'd245;
     memory[1254] = 32'd53;
     memory[1255] = 32'd216;
     memory[1256] = 32'd184;
     memory[1257] = 32'd188;
     memory[1258] = 32'd253;
     memory[1259] = 32'd148;
     memory[1260] = 32'd180;
     memory[1261] = 32'd50;
     memory[1262] = 32'd151;
     memory[1263] = 32'd254;
     memory[1264] = 32'd143;
     memory[1265] = 32'd209;
     memory[1266] = 32'd74;
     memory[1267] = 32'd205;
     memory[1268] = 32'd120;
     memory[1269] = 32'd235;
     memory[1270] = 32'd245;
     memory[1271] = 32'd200;
     memory[1272] = 32'd23;
     memory[1273] = 32'd198;
     memory[1274] = 32'd125;
     memory[1275] = 32'd118;
     memory[1276] = 32'd222;
     memory[1277] = 32'd235;
     memory[1278] = 32'd104;
     memory[1279] = 32'd47;
     memory[1280] = 32'd51;
     memory[1281] = 32'd10;
     memory[1282] = 32'd72;
     memory[1283] = 32'd33;
     memory[1284] = 32'd100;
     memory[1285] = 32'd191;
     memory[1286] = 32'd170;
     memory[1287] = 32'd20;
     memory[1288] = 32'd33;
     memory[1289] = 32'd91;
     memory[1290] = 32'd32;
     memory[1291] = 32'd128;
     memory[1292] = 32'd56;
     memory[1293] = 32'd150;
     memory[1294] = 32'd202;
     memory[1295] = 32'd87;
     memory[1296] = 32'd43;
     memory[1297] = 32'd214;
     memory[1298] = 32'd147;
     memory[1299] = 32'd192;
     memory[1300] = 32'd204;
     memory[1301] = 32'd69;
     memory[1302] = 32'd26;
     memory[1303] = 32'd72;
     memory[1304] = 32'd249;
     memory[1305] = 32'd180;
     memory[1306] = 32'd248;
     memory[1307] = 32'd41;
     memory[1308] = 32'd125;
     memory[1309] = 32'd50;
     memory[1310] = 32'd175;
     memory[1311] = 32'd166;
     memory[1312] = 32'd127;
     memory[1313] = 32'd114;
     memory[1314] = 32'd229;
     memory[1315] = 32'd254;
     memory[1316] = 32'd167;
     memory[1317] = 32'd162;
     memory[1318] = 32'd252;
     memory[1319] = 32'd136;
     memory[1320] = 32'd8;
     memory[1321] = 32'd3;
     memory[1322] = 32'd44;
     memory[1323] = 32'd112;
     memory[1324] = 32'd77;
     memory[1325] = 32'd232;
     memory[1326] = 32'd247;
     memory[1327] = 32'd84;
     memory[1328] = 32'd46;
     memory[1329] = 32'd34;
     memory[1330] = 32'd61;
     memory[1331] = 32'd233;
     memory[1332] = 32'd126;
     memory[1333] = 32'd34;
     memory[1334] = 32'd136;
     memory[1335] = 32'd43;
     memory[1336] = 32'd96;
     memory[1337] = 32'd15;
     memory[1338] = 32'd173;
     memory[1339] = 32'd120;
     memory[1340] = 32'd79;
     memory[1341] = 32'd120;
     memory[1342] = 32'd130;
     memory[1343] = 32'd110;
     memory[1344] = 32'd254;
     memory[1345] = 32'd8;
     memory[1346] = 32'd121;
     memory[1347] = 32'd153;
     memory[1348] = 32'd211;
     memory[1349] = 32'd176;
     memory[1350] = 32'd82;
     memory[1351] = 32'd171;
     memory[1352] = 32'd209;
     memory[1353] = 32'd142;
     memory[1354] = 32'd156;
     memory[1355] = 32'd218;
     memory[1356] = 32'd169;
     memory[1357] = 32'd77;
     memory[1358] = 32'd195;
     memory[1359] = 32'd210;
     memory[1360] = 32'd14;
     memory[1361] = 32'd99;
     memory[1362] = 32'd130;
     memory[1363] = 32'd178;
     memory[1364] = 32'd140;
     memory[1365] = 32'd171;
     memory[1366] = 32'd56;
     memory[1367] = 32'd41;
     memory[1368] = 32'd38;
     memory[1369] = 32'd64;
     memory[1370] = 32'd73;
     memory[1371] = 32'd97;
     memory[1372] = 32'd136;
     memory[1373] = 32'd120;
     memory[1374] = 32'd8;
     memory[1375] = 32'd142;
     memory[1376] = 32'd159;
     memory[1377] = 32'd234;
     memory[1378] = 32'd116;
     memory[1379] = 32'd154;
     memory[1380] = 32'd231;
     memory[1381] = 32'd13;
     memory[1382] = 32'd17;
     memory[1383] = 32'd91;
     memory[1384] = 32'd49;
     memory[1385] = 32'd209;
     memory[1386] = 32'd16;
     memory[1387] = 32'd7;
     memory[1388] = 32'd61;
     memory[1389] = 32'd233;
     memory[1390] = 32'd222;
     memory[1391] = 32'd187;
     memory[1392] = 32'd60;
     memory[1393] = 32'd55;
     memory[1394] = 32'd50;
     memory[1395] = 32'd153;
     memory[1396] = 32'd238;
     memory[1397] = 32'd193;
     memory[1398] = 32'd37;
     memory[1399] = 32'd225;
     memory[1400] = 32'd122;
     memory[1401] = 32'd144;
     memory[1402] = 32'd161;
     memory[1403] = 32'd41;
     memory[1404] = 32'd27;
     memory[1405] = 32'd59;
     memory[1406] = 32'd156;
     memory[1407] = 32'd18;
     memory[1408] = 32'd149;
     memory[1409] = 32'd115;
     memory[1410] = 32'd188;
     memory[1411] = 32'd25;
     memory[1412] = 32'd136;
     memory[1413] = 32'd233;
     memory[1414] = 32'd98;
     memory[1415] = 32'd152;
     memory[1416] = 32'd133;
     memory[1417] = 32'd23;
     memory[1418] = 32'd198;
     memory[1419] = 32'd75;
     memory[1420] = 32'd242;
     memory[1421] = 32'd188;
     memory[1422] = 32'd74;
     memory[1423] = 32'd154;
     memory[1424] = 32'd16;
     memory[1425] = 32'd71;
     memory[1426] = 32'd164;
     memory[1427] = 32'd236;
     memory[1428] = 32'd187;
     memory[1429] = 32'd254;
     memory[1430] = 32'd2;
     memory[1431] = 32'd50;
     memory[1432] = 32'd174;
     memory[1433] = 32'd206;
     memory[1434] = 32'd100;
     memory[1435] = 32'd119;
     memory[1436] = 32'd196;
     memory[1437] = 32'd178;
     memory[1438] = 32'd176;
     memory[1439] = 32'd227;
     memory[1440] = 32'd166;
     memory[1441] = 32'd183;
     memory[1442] = 32'd132;
     memory[1443] = 32'd192;
     memory[1444] = 32'd94;
     memory[1445] = 32'd214;
     memory[1446] = 32'd74;
     memory[1447] = 32'd175;
     memory[1448] = 32'd198;
     memory[1449] = 32'd183;
     memory[1450] = 32'd36;
     memory[1451] = 32'd222;
     memory[1452] = 32'd214;
     memory[1453] = 32'd0;
     memory[1454] = 32'd239;
     memory[1455] = 32'd107;
     memory[1456] = 32'd212;
     memory[1457] = 32'd114;
     memory[1458] = 32'd111;
     memory[1459] = 32'd130;
     memory[1460] = 32'd136;
     memory[1461] = 32'd222;
     memory[1462] = 32'd213;
     memory[1463] = 32'd85;
     memory[1464] = 32'd115;
     memory[1465] = 32'd11;
     memory[1466] = 32'd99;
     memory[1467] = 32'd69;
     memory[1468] = 32'd232;
     memory[1469] = 32'd228;
     memory[1470] = 32'd18;
     memory[1471] = 32'd37;
     memory[1472] = 32'd76;
     memory[1473] = 32'd81;
     memory[1474] = 32'd126;
     memory[1475] = 32'd74;
     memory[1476] = 32'd215;
     memory[1477] = 32'd181;
     memory[1478] = 32'd53;
     memory[1479] = 32'd111;
     memory[1480] = 32'd156;
     memory[1481] = 32'd140;
     memory[1482] = 32'd14;
     memory[1483] = 32'd136;
     memory[1484] = 32'd134;
     memory[1485] = 32'd56;
     memory[1486] = 32'd93;
     memory[1487] = 32'd65;
     memory[1488] = 32'd102;
     memory[1489] = 32'd207;
     memory[1490] = 32'd65;
     memory[1491] = 32'd100;
     memory[1492] = 32'd93;
     memory[1493] = 32'd28;
     memory[1494] = 32'd150;
     memory[1495] = 32'd238;
     memory[1496] = 32'd28;
     memory[1497] = 32'd13;
     memory[1498] = 32'd48;
     memory[1499] = 32'd254;
     memory[1500] = 32'd247;
     memory[1501] = 32'd116;
     memory[1502] = 32'd158;
     memory[1503] = 32'd128;
     memory[1504] = 32'd45;
     memory[1505] = 32'd190;
     memory[1506] = 32'd164;
     memory[1507] = 32'd171;
     memory[1508] = 32'd211;
     memory[1509] = 32'd176;
     memory[1510] = 32'd178;
     memory[1511] = 32'd182;
     memory[1512] = 32'd29;
     memory[1513] = 32'd204;
     memory[1514] = 32'd229;
     memory[1515] = 32'd31;
     memory[1516] = 32'd147;
     memory[1517] = 32'd245;
     memory[1518] = 32'd137;
     memory[1519] = 32'd118;
     memory[1520] = 32'd5;
     memory[1521] = 32'd163;
     memory[1522] = 32'd117;
     memory[1523] = 32'd196;
     memory[1524] = 32'd57;
     memory[1525] = 32'd183;
     memory[1526] = 32'd184;
     memory[1527] = 32'd47;
     memory[1528] = 32'd67;
     memory[1529] = 32'd247;
     memory[1530] = 32'd201;
     memory[1531] = 32'd38;
     memory[1532] = 32'd92;
     memory[1533] = 32'd11;
     memory[1534] = 32'd123;
     memory[1535] = 32'd114;
     memory[1536] = 32'd49;
     memory[1537] = 32'd1;
     memory[1538] = 32'd231;
     memory[1539] = 32'd131;
     memory[1540] = 32'd229;
     memory[1541] = 32'd219;
     memory[1542] = 32'd115;
     memory[1543] = 32'd104;
     memory[1544] = 32'd3;
     memory[1545] = 32'd179;
     memory[1546] = 32'd136;
     memory[1547] = 32'd236;
     memory[1548] = 32'd197;
     memory[1549] = 32'd70;
     memory[1550] = 32'd120;
     memory[1551] = 32'd227;
     memory[1552] = 32'd147;
     memory[1553] = 32'd121;
     memory[1554] = 32'd142;
     memory[1555] = 32'd84;
     memory[1556] = 32'd146;
     memory[1557] = 32'd113;
     memory[1558] = 32'd243;
     memory[1559] = 32'd81;
     memory[1560] = 32'd204;
     memory[1561] = 32'd73;
     memory[1562] = 32'd214;
     memory[1563] = 32'd121;
     memory[1564] = 32'd169;
     memory[1565] = 32'd191;
     memory[1566] = 32'd35;
     memory[1567] = 32'd113;
     memory[1568] = 32'd248;
     memory[1569] = 32'd78;
     memory[1570] = 32'd69;
     memory[1571] = 32'd56;
     memory[1572] = 32'd17;
     memory[1573] = 32'd40;
     memory[1574] = 32'd147;
     memory[1575] = 32'd177;
     memory[1576] = 32'd96;
     memory[1577] = 32'd206;
     memory[1578] = 32'd160;
     memory[1579] = 32'd116;
     memory[1580] = 32'd199;
     memory[1581] = 32'd53;
     memory[1582] = 32'd192;
     memory[1583] = 32'd88;
     memory[1584] = 32'd188;
     memory[1585] = 32'd65;
     memory[1586] = 32'd102;
     memory[1587] = 32'd23;
     memory[1588] = 32'd55;
     memory[1589] = 32'd191;
     memory[1590] = 32'd45;
     memory[1591] = 32'd39;
     memory[1592] = 32'd88;
     memory[1593] = 32'd238;
     memory[1594] = 32'd205;
     memory[1595] = 32'd84;
     memory[1596] = 32'd210;
     memory[1597] = 32'd179;
     memory[1598] = 32'd49;
     memory[1599] = 32'd176;
     memory[1600] = 32'd52;
     memory[1601] = 32'd162;
     memory[1602] = 32'd48;
     memory[1603] = 32'd227;
     memory[1604] = 32'd132;
     memory[1605] = 32'd192;
     memory[1606] = 32'd94;
     memory[1607] = 32'd243;
     memory[1608] = 32'd44;
     memory[1609] = 32'd140;
     memory[1610] = 32'd34;
     memory[1611] = 32'd196;
     memory[1612] = 32'd106;
     memory[1613] = 32'd182;
     memory[1614] = 32'd38;
     memory[1615] = 32'd4;
     memory[1616] = 32'd58;
     memory[1617] = 32'd129;
     memory[1618] = 32'd240;
     memory[1619] = 32'd173;
     memory[1620] = 32'd121;
     memory[1621] = 32'd109;
     memory[1622] = 32'd205;
     memory[1623] = 32'd112;
     memory[1624] = 32'd13;
     memory[1625] = 32'd163;
     memory[1626] = 32'd153;
     memory[1627] = 32'd24;
     memory[1628] = 32'd230;
     memory[1629] = 32'd20;
     memory[1630] = 32'd253;
     memory[1631] = 32'd49;
     memory[1632] = 32'd184;
     memory[1633] = 32'd14;
     memory[1634] = 32'd10;
     memory[1635] = 32'd96;
     memory[1636] = 32'd94;
     memory[1637] = 32'd178;
     memory[1638] = 32'd159;
     memory[1639] = 32'd80;
     memory[1640] = 32'd146;
     memory[1641] = 32'd91;
     memory[1642] = 32'd171;
     memory[1643] = 32'd235;
     memory[1644] = 32'd20;
     memory[1645] = 32'd150;
     memory[1646] = 32'd135;
     memory[1647] = 32'd41;
     memory[1648] = 32'd155;
     memory[1649] = 32'd93;
     memory[1650] = 32'd120;
     memory[1651] = 32'd184;
     memory[1652] = 32'd172;
     memory[1653] = 32'd55;
     memory[1654] = 32'd113;
     memory[1655] = 32'd47;
     memory[1656] = 32'd99;
     memory[1657] = 32'd70;
     memory[1658] = 32'd208;
     memory[1659] = 32'd71;
     memory[1660] = 32'd188;
     memory[1661] = 32'd92;
     memory[1662] = 32'd208;
     memory[1663] = 32'd247;
     memory[1664] = 32'd96;
     memory[1665] = 32'd81;
     memory[1666] = 32'd12;
     memory[1667] = 32'd5;
     memory[1668] = 32'd64;
     memory[1669] = 32'd70;
     memory[1670] = 32'd209;
     memory[1671] = 32'd146;
     memory[1672] = 32'd185;
     memory[1673] = 32'd142;
     memory[1674] = 32'd25;
     memory[1675] = 32'd198;
     memory[1676] = 32'd16;
     memory[1677] = 32'd64;
     memory[1678] = 32'd92;
     memory[1679] = 32'd152;
     memory[1680] = 32'd144;
     memory[1681] = 32'd26;
     memory[1682] = 32'd243;
     memory[1683] = 32'd9;
     memory[1684] = 32'd21;
     memory[1685] = 32'd73;
     memory[1686] = 32'd113;
     memory[1687] = 32'd171;
     memory[1688] = 32'd32;
     memory[1689] = 32'd149;
     memory[1690] = 32'd110;
     memory[1691] = 32'd170;
     memory[1692] = 32'd33;
     memory[1693] = 32'd128;
     memory[1694] = 32'd232;
     memory[1695] = 32'd132;
     memory[1696] = 32'd42;
     memory[1697] = 32'd206;
     memory[1698] = 32'd174;
     memory[1699] = 32'd249;
     memory[1700] = 32'd126;
     memory[1701] = 32'd222;
     memory[1702] = 32'd108;
     memory[1703] = 32'd106;
     memory[1704] = 32'd38;
     memory[1705] = 32'd78;
     memory[1706] = 32'd163;
     memory[1707] = 32'd181;
     memory[1708] = 32'd69;
     memory[1709] = 32'd60;
     memory[1710] = 32'd203;
     memory[1711] = 32'd94;
     memory[1712] = 32'd118;
     memory[1713] = 32'd252;
     memory[1714] = 32'd135;
     memory[1715] = 32'd45;
     memory[1716] = 32'd123;
     memory[1717] = 32'd148;
     memory[1718] = 32'd27;
     memory[1719] = 32'd37;
     memory[1720] = 32'd232;
     memory[1721] = 32'd36;
     memory[1722] = 32'd122;
     memory[1723] = 32'd30;
     memory[1724] = 32'd207;
     memory[1725] = 32'd146;
     memory[1726] = 32'd224;
     memory[1727] = 32'd156;
     memory[1728] = 32'd183;
     memory[1729] = 32'd19;
     memory[1730] = 32'd38;
     memory[1731] = 32'd105;
     memory[1732] = 32'd174;
     memory[1733] = 32'd113;
     memory[1734] = 32'd58;
     memory[1735] = 32'd209;
     memory[1736] = 32'd40;
     memory[1737] = 32'd253;
     memory[1738] = 32'd73;
     memory[1739] = 32'd229;
     memory[1740] = 32'd20;
     memory[1741] = 32'd154;
     memory[1742] = 32'd81;
     memory[1743] = 32'd139;
     memory[1744] = 32'd55;
     memory[1745] = 32'd87;
     memory[1746] = 32'd144;
     memory[1747] = 32'd109;
     memory[1748] = 32'd95;
     memory[1749] = 32'd51;
     memory[1750] = 32'd74;
     memory[1751] = 32'd171;
     memory[1752] = 32'd106;
     memory[1753] = 32'd95;
     memory[1754] = 32'd146;
     memory[1755] = 32'd207;
     memory[1756] = 32'd98;
     memory[1757] = 32'd106;
     memory[1758] = 32'd178;
     memory[1759] = 32'd199;
     memory[1760] = 32'd135;
     memory[1761] = 32'd56;
     memory[1762] = 32'd108;
     memory[1763] = 32'd186;
     memory[1764] = 32'd186;
     memory[1765] = 32'd167;
     memory[1766] = 32'd249;
     memory[1767] = 32'd244;
     memory[1768] = 32'd204;
     memory[1769] = 32'd62;
     memory[1770] = 32'd222;
     memory[1771] = 32'd205;
     memory[1772] = 32'd94;
     memory[1773] = 32'd11;
     memory[1774] = 32'd245;
     memory[1775] = 32'd202;
     memory[1776] = 32'd238;
     memory[1777] = 32'd141;
     memory[1778] = 32'd220;
     memory[1779] = 32'd92;
     memory[1780] = 32'd190;
     memory[1781] = 32'd155;
     memory[1782] = 32'd218;
     memory[1783] = 32'd201;
     memory[1784] = 32'd128;
     memory[1785] = 32'd240;
     memory[1786] = 32'd47;
     memory[1787] = 32'd150;
     memory[1788] = 32'd90;
     memory[1789] = 32'd55;
     memory[1790] = 32'd108;
     memory[1791] = 32'd244;
     memory[1792] = 32'd190;
     memory[1793] = 32'd119;
     memory[1794] = 32'd17;
     memory[1795] = 32'd25;
     memory[1796] = 32'd175;
     memory[1797] = 32'd250;
     memory[1798] = 32'd169;
     memory[1799] = 32'd207;
     memory[1800] = 32'd6;
     memory[1801] = 32'd168;
     memory[1802] = 32'd194;
     memory[1803] = 32'd171;
     memory[1804] = 32'd159;
     memory[1805] = 32'd182;
     memory[1806] = 32'd17;
     memory[1807] = 32'd2;
     memory[1808] = 32'd38;
     memory[1809] = 32'd227;
     memory[1810] = 32'd18;
     memory[1811] = 32'd132;
     memory[1812] = 32'd198;
     memory[1813] = 32'd244;
     memory[1814] = 32'd192;
     memory[1815] = 32'd187;
     memory[1816] = 32'd89;
     memory[1817] = 32'd232;
     memory[1818] = 32'd97;
     memory[1819] = 32'd46;
     memory[1820] = 32'd19;
     memory[1821] = 32'd66;
     memory[1822] = 32'd33;
     memory[1823] = 32'd231;
     memory[1824] = 32'd188;
     memory[1825] = 32'd80;
     memory[1826] = 32'd34;
     memory[1827] = 32'd196;
     memory[1828] = 32'd7;
     memory[1829] = 32'd14;
     memory[1830] = 32'd203;
     memory[1831] = 32'd93;
     memory[1832] = 32'd229;
     memory[1833] = 32'd75;
     memory[1834] = 32'd97;
     memory[1835] = 32'd44;
     memory[1836] = 32'd214;
     memory[1837] = 32'd243;
     memory[1838] = 32'd101;
     memory[1839] = 32'd118;
     memory[1840] = 32'd212;
     memory[1841] = 32'd237;
     memory[1842] = 32'd161;
     memory[1843] = 32'd253;
     memory[1844] = 32'd165;
     memory[1845] = 32'd230;
     memory[1846] = 32'd13;
     memory[1847] = 32'd229;
     memory[1848] = 32'd199;
     memory[1849] = 32'd221;
     memory[1850] = 32'd151;
     memory[1851] = 32'd181;
     memory[1852] = 32'd94;
     memory[1853] = 32'd163;
     memory[1854] = 32'd82;
     memory[1855] = 32'd226;
     memory[1856] = 32'd248;
     memory[1857] = 32'd32;
     memory[1858] = 32'd127;
     memory[1859] = 32'd138;
     memory[1860] = 32'd202;
     memory[1861] = 32'd161;
     memory[1862] = 32'd69;
     memory[1863] = 32'd55;
     memory[1864] = 32'd50;
     memory[1865] = 32'd188;
     memory[1866] = 32'd135;
     memory[1867] = 32'd98;
     memory[1868] = 32'd4;
     memory[1869] = 32'd224;
     memory[1870] = 32'd190;
     memory[1871] = 32'd237;
     memory[1872] = 32'd218;
     memory[1873] = 32'd113;
     memory[1874] = 32'd239;
     memory[1875] = 32'd53;
     memory[1876] = 32'd175;
     memory[1877] = 32'd53;
     memory[1878] = 32'd162;
     memory[1879] = 32'd243;
     memory[1880] = 32'd79;
     memory[1881] = 32'd154;
     memory[1882] = 32'd70;
     memory[1883] = 32'd222;
     memory[1884] = 32'd221;
     memory[1885] = 32'd186;
     memory[1886] = 32'd98;
     memory[1887] = 32'd13;
     memory[1888] = 32'd32;
     memory[1889] = 32'd165;
     memory[1890] = 32'd231;
     memory[1891] = 32'd217;
     memory[1892] = 32'd11;
     memory[1893] = 32'd186;
     memory[1894] = 32'd154;
     memory[1895] = 32'd190;
     memory[1896] = 32'd209;
     memory[1897] = 32'd164;
     memory[1898] = 32'd242;
     memory[1899] = 32'd134;
     memory[1900] = 32'd175;
     memory[1901] = 32'd93;
     memory[1902] = 32'd19;
     memory[1903] = 32'd227;
     memory[1904] = 32'd48;
     memory[1905] = 32'd37;
     memory[1906] = 32'd214;
     memory[1907] = 32'd254;
     memory[1908] = 32'd83;
     memory[1909] = 32'd193;
     memory[1910] = 32'd63;
     memory[1911] = 32'd199;
     memory[1912] = 32'd105;
     memory[1913] = 32'd248;
     memory[1914] = 32'd190;
     memory[1915] = 32'd117;
     memory[1916] = 32'd214;
     memory[1917] = 32'd111;
     memory[1918] = 32'd6;
     memory[1919] = 32'd47;
     memory[1920] = 32'd14;
     memory[1921] = 32'd217;
     memory[1922] = 32'd79;
     memory[1923] = 32'd197;
     memory[1924] = 32'd39;
     memory[1925] = 32'd239;
     memory[1926] = 32'd212;
     memory[1927] = 32'd201;
     memory[1928] = 32'd73;
     memory[1929] = 32'd128;
     memory[1930] = 32'd248;
     memory[1931] = 32'd211;
     memory[1932] = 32'd210;
     memory[1933] = 32'd207;
     memory[1934] = 32'd105;
     memory[1935] = 32'd166;
     memory[1936] = 32'd103;
     memory[1937] = 32'd192;
     memory[1938] = 32'd186;
     memory[1939] = 32'd163;
     memory[1940] = 32'd94;
     memory[1941] = 32'd153;
     memory[1942] = 32'd231;
     memory[1943] = 32'd3;
     memory[1944] = 32'd127;
     memory[1945] = 32'd168;
     memory[1946] = 32'd97;
     memory[1947] = 32'd74;
     memory[1948] = 32'd177;
     memory[1949] = 32'd142;
     memory[1950] = 32'd126;
     memory[1951] = 32'd245;
     memory[1952] = 32'd37;
     memory[1953] = 32'd101;
     memory[1954] = 32'd215;
     memory[1955] = 32'd72;
     memory[1956] = 32'd4;
     memory[1957] = 32'd180;
     memory[1958] = 32'd23;
     memory[1959] = 32'd28;
     memory[1960] = 32'd173;
     memory[1961] = 32'd141;
     memory[1962] = 32'd185;
     memory[1963] = 32'd39;
     memory[1964] = 32'd97;
     memory[1965] = 32'd64;
     memory[1966] = 32'd53;
     memory[1967] = 32'd187;
     memory[1968] = 32'd18;
     memory[1969] = 32'd229;
     memory[1970] = 32'd92;
     memory[1971] = 32'd155;
     memory[1972] = 32'd55;
     memory[1973] = 32'd228;
     memory[1974] = 32'd188;
     memory[1975] = 32'd129;
     memory[1976] = 32'd109;
     memory[1977] = 32'd134;
     memory[1978] = 32'd36;
     memory[1979] = 32'd192;
     memory[1980] = 32'd248;
     memory[1981] = 32'd153;
     memory[1982] = 32'd204;
     memory[1983] = 32'd81;
     memory[1984] = 32'd3;
     memory[1985] = 32'd183;
     memory[1986] = 32'd57;
     memory[1987] = 32'd215;
     memory[1988] = 32'd83;
     memory[1989] = 32'd215;
     memory[1990] = 32'd28;
     memory[1991] = 32'd99;
     memory[1992] = 32'd54;
     memory[1993] = 32'd15;
     memory[1994] = 32'd254;
     memory[1995] = 32'd30;
     memory[1996] = 32'd113;
     memory[1997] = 32'd224;
     memory[1998] = 32'd25;
     memory[1999] = 32'd96;
     memory[2000] = 32'd10;
     memory[2001] = 32'd84;
     memory[2002] = 32'd250;
     memory[2003] = 32'd114;
     memory[2004] = 32'd26;
     memory[2005] = 32'd29;
     memory[2006] = 32'd89;
     memory[2007] = 32'd139;
     memory[2008] = 32'd133;
     memory[2009] = 32'd125;
     memory[2010] = 32'd43;
     memory[2011] = 32'd129;
     memory[2012] = 32'd212;
     memory[2013] = 32'd223;
     memory[2014] = 32'd51;
     memory[2015] = 32'd61;
     memory[2016] = 32'd99;
     memory[2017] = 32'd58;
     memory[2018] = 32'd72;
     memory[2019] = 32'd146;
     memory[2020] = 32'd0;
     memory[2021] = 32'd200;
     memory[2022] = 32'd160;
     memory[2023] = 32'd189;
     memory[2024] = 32'd94;
     memory[2025] = 32'd149;
     memory[2026] = 32'd142;
     memory[2027] = 32'd54;
     memory[2028] = 32'd202;
     memory[2029] = 32'd0;
     memory[2030] = 32'd201;
     memory[2031] = 32'd133;
     memory[2032] = 32'd68;
     memory[2033] = 32'd30;
     memory[2034] = 32'd110;
     memory[2035] = 32'd38;
     memory[2036] = 32'd127;
     memory[2037] = 32'd169;
     memory[2038] = 32'd253;
     memory[2039] = 32'd159;
     memory[2040] = 32'd144;
     memory[2041] = 32'd193;
     memory[2042] = 32'd210;
     memory[2043] = 32'd222;
     memory[2044] = 32'd200;
     memory[2045] = 32'd32;
     memory[2046] = 32'd245;
     memory[2047] = 32'd35;
     memory[2048] = 32'd240;
     memory[2049] = 32'd229;
     memory[2050] = 32'd201;
     memory[2051] = 32'd102;
     memory[2052] = 32'd66;
     memory[2053] = 32'd23;
     memory[2054] = 32'd243;
     memory[2055] = 32'd167;
     memory[2056] = 32'd67;
     memory[2057] = 32'd143;
     memory[2058] = 32'd31;
     memory[2059] = 32'd231;
     memory[2060] = 32'd101;
     memory[2061] = 32'd203;
     memory[2062] = 32'd149;
     memory[2063] = 32'd14;
     memory[2064] = 32'd106;
     memory[2065] = 32'd76;
     memory[2066] = 32'd102;
     memory[2067] = 32'd249;
     memory[2068] = 32'd180;
     memory[2069] = 32'd175;
     memory[2070] = 32'd225;
     memory[2071] = 32'd89;
     memory[2072] = 32'd152;
     memory[2073] = 32'd205;
     memory[2074] = 32'd172;
     memory[2075] = 32'd119;
     memory[2076] = 32'd0;
     memory[2077] = 32'd51;
     memory[2078] = 32'd8;
     memory[2079] = 32'd91;
     memory[2080] = 32'd48;
     memory[2081] = 32'd19;
     memory[2082] = 32'd87;
     memory[2083] = 32'd150;
     memory[2084] = 32'd226;
     memory[2085] = 32'd253;
     memory[2086] = 32'd217;
     memory[2087] = 32'd158;
     memory[2088] = 32'd175;
     memory[2089] = 32'd231;
     memory[2090] = 32'd23;
     memory[2091] = 32'd107;
     memory[2092] = 32'd164;
     memory[2093] = 32'd233;
     memory[2094] = 32'd171;
     memory[2095] = 32'd114;
     memory[2096] = 32'd135;
     memory[2097] = 32'd53;
     memory[2098] = 32'd229;
     memory[2099] = 32'd126;
     memory[2100] = 32'd181;
     memory[2101] = 32'd108;
     memory[2102] = 32'd117;
     memory[2103] = 32'd187;
     memory[2104] = 32'd241;
     memory[2105] = 32'd225;
     memory[2106] = 32'd110;
     memory[2107] = 32'd72;
     memory[2108] = 32'd109;
     memory[2109] = 32'd47;
     memory[2110] = 32'd15;
     memory[2111] = 32'd153;
     memory[2112] = 32'd214;
     memory[2113] = 32'd15;
     memory[2114] = 32'd57;
     memory[2115] = 32'd139;
     memory[2116] = 32'd196;
     memory[2117] = 32'd115;
     memory[2118] = 32'd142;
     memory[2119] = 32'd166;
     memory[2120] = 32'd207;
     memory[2121] = 32'd175;
     memory[2122] = 32'd252;
     memory[2123] = 32'd72;
     memory[2124] = 32'd0;
     memory[2125] = 32'd83;
     memory[2126] = 32'd162;
     memory[2127] = 32'd169;
     memory[2128] = 32'd96;
     memory[2129] = 32'd171;
     memory[2130] = 32'd11;
     memory[2131] = 32'd48;
     memory[2132] = 32'd198;
     memory[2133] = 32'd122;
     memory[2134] = 32'd19;
     memory[2135] = 32'd50;
     memory[2136] = 32'd170;
     memory[2137] = 32'd116;
     memory[2138] = 32'd252;
     memory[2139] = 32'd236;
     memory[2140] = 32'd108;
     memory[2141] = 32'd187;
     memory[2142] = 32'd248;
     memory[2143] = 32'd253;
     memory[2144] = 32'd115;
     memory[2145] = 32'd55;
     memory[2146] = 32'd170;
     memory[2147] = 32'd252;
     memory[2148] = 32'd20;
     memory[2149] = 32'd240;
     memory[2150] = 32'd4;
     memory[2151] = 32'd199;
     memory[2152] = 32'd229;
     memory[2153] = 32'd157;
     memory[2154] = 32'd190;
     memory[2155] = 32'd203;
     memory[2156] = 32'd166;
     memory[2157] = 32'd45;
     memory[2158] = 32'd46;
     memory[2159] = 32'd173;
     memory[2160] = 32'd17;
     memory[2161] = 32'd83;
     memory[2162] = 32'd88;
     memory[2163] = 32'd217;
     memory[2164] = 32'd63;
     memory[2165] = 32'd21;
     memory[2166] = 32'd133;
     memory[2167] = 32'd193;
     memory[2168] = 32'd222;
     memory[2169] = 32'd114;
     memory[2170] = 32'd69;
     memory[2171] = 32'd37;
     memory[2172] = 32'd193;
     memory[2173] = 32'd197;
     memory[2174] = 32'd215;
     memory[2175] = 32'd154;
     memory[2176] = 32'd99;
     memory[2177] = 32'd218;
     memory[2178] = 32'd252;
     memory[2179] = 32'd76;
     memory[2180] = 32'd245;
     memory[2181] = 32'd36;
     memory[2182] = 32'd67;
     memory[2183] = 32'd102;
     memory[2184] = 32'd166;
     memory[2185] = 32'd67;
     memory[2186] = 32'd20;
     memory[2187] = 32'd236;
     memory[2188] = 32'd48;
     memory[2189] = 32'd252;
     memory[2190] = 32'd223;
     memory[2191] = 32'd140;
     memory[2192] = 32'd81;
     memory[2193] = 32'd148;
     memory[2194] = 32'd16;
     memory[2195] = 32'd116;
     memory[2196] = 32'd72;
     memory[2197] = 32'd154;
     memory[2198] = 32'd251;
     memory[2199] = 32'd71;
     memory[2200] = 32'd229;
     memory[2201] = 32'd6;
     memory[2202] = 32'd120;
     memory[2203] = 32'd22;
     memory[2204] = 32'd194;
     memory[2205] = 32'd172;
     memory[2206] = 32'd72;
     memory[2207] = 32'd58;
     memory[2208] = 32'd7;
     memory[2209] = 32'd118;
     memory[2210] = 32'd139;
     memory[2211] = 32'd176;
     memory[2212] = 32'd209;
     memory[2213] = 32'd131;
     memory[2214] = 32'd72;
     memory[2215] = 32'd95;
     memory[2216] = 32'd43;
     memory[2217] = 32'd168;
     memory[2218] = 32'd19;
     memory[2219] = 32'd205;
     memory[2220] = 32'd224;
     memory[2221] = 32'd242;
     memory[2222] = 32'd209;
     memory[2223] = 32'd130;
     memory[2224] = 32'd217;
     memory[2225] = 32'd173;
     memory[2226] = 32'd22;
     memory[2227] = 32'd80;
     memory[2228] = 32'd7;
     memory[2229] = 32'd74;
     memory[2230] = 32'd73;
     memory[2231] = 32'd96;
     memory[2232] = 32'd123;
     memory[2233] = 32'd159;
     memory[2234] = 32'd94;
     memory[2235] = 32'd55;
     memory[2236] = 32'd115;
     memory[2237] = 32'd194;
     memory[2238] = 32'd27;
     memory[2239] = 32'd182;
     memory[2240] = 32'd95;
     memory[2241] = 32'd181;
     memory[2242] = 32'd167;
     memory[2243] = 32'd38;
     memory[2244] = 32'd232;
     memory[2245] = 32'd84;
     memory[2246] = 32'd136;
     memory[2247] = 32'd169;
     memory[2248] = 32'd224;
     memory[2249] = 32'd167;
     memory[2250] = 32'd240;
     memory[2251] = 32'd131;
     memory[2252] = 32'd153;
     memory[2253] = 32'd213;
     memory[2254] = 32'd132;
     memory[2255] = 32'd203;
     memory[2256] = 32'd191;
     memory[2257] = 32'd216;
     memory[2258] = 32'd203;
     memory[2259] = 32'd150;
     memory[2260] = 32'd209;
     memory[2261] = 32'd60;
     memory[2262] = 32'd170;
     memory[2263] = 32'd205;
     memory[2264] = 32'd240;
     memory[2265] = 32'd149;
     memory[2266] = 32'd85;
     memory[2267] = 32'd192;
     memory[2268] = 32'd55;
     memory[2269] = 32'd154;
     memory[2270] = 32'd14;
     memory[2271] = 32'd6;
     memory[2272] = 32'd219;
     memory[2273] = 32'd187;
     memory[2274] = 32'd5;
     memory[2275] = 32'd11;
     memory[2276] = 32'd235;
     memory[2277] = 32'd45;
     memory[2278] = 32'd154;
     memory[2279] = 32'd30;
     memory[2280] = 32'd76;
     memory[2281] = 32'd106;
     memory[2282] = 32'd16;
     memory[2283] = 32'd213;
     memory[2284] = 32'd193;
     memory[2285] = 32'd90;
     memory[2286] = 32'd102;
     memory[2287] = 32'd79;
     memory[2288] = 32'd126;
     memory[2289] = 32'd46;
     memory[2290] = 32'd212;
     memory[2291] = 32'd16;
     memory[2292] = 32'd94;
     memory[2293] = 32'd51;
     memory[2294] = 32'd225;
     memory[2295] = 32'd122;
     memory[2296] = 32'd192;
     memory[2297] = 32'd123;
     memory[2298] = 32'd56;
     memory[2299] = 32'd239;
     memory[2300] = 32'd65;
     memory[2301] = 32'd218;
     memory[2302] = 32'd158;
     memory[2303] = 32'd168;
     memory[2304] = 32'd246;
     memory[2305] = 32'd20;
     memory[2306] = 32'd21;
     memory[2307] = 32'd211;
     memory[2308] = 32'd67;
     memory[2309] = 32'd111;
     memory[2310] = 32'd133;
     memory[2311] = 32'd224;
     memory[2312] = 32'd49;
     memory[2313] = 32'd250;
     memory[2314] = 32'd198;
     memory[2315] = 32'd115;
     memory[2316] = 32'd53;
     memory[2317] = 32'd142;
     memory[2318] = 32'd92;
     memory[2319] = 32'd56;
     memory[2320] = 32'd81;
     memory[2321] = 32'd76;
     memory[2322] = 32'd49;
     memory[2323] = 32'd252;
     memory[2324] = 32'd117;
     memory[2325] = 32'd42;
     memory[2326] = 32'd248;
     memory[2327] = 32'd167;
     memory[2328] = 32'd213;
     memory[2329] = 32'd35;
     memory[2330] = 32'd73;
     memory[2331] = 32'd228;
     memory[2332] = 32'd154;
     memory[2333] = 32'd245;
     memory[2334] = 32'd116;
     memory[2335] = 32'd65;
     memory[2336] = 32'd115;
     memory[2337] = 32'd54;
     memory[2338] = 32'd186;
     memory[2339] = 32'd68;
     memory[2340] = 32'd59;
     memory[2341] = 32'd163;
     memory[2342] = 32'd117;
     memory[2343] = 32'd66;
     memory[2344] = 32'd148;
     memory[2345] = 32'd235;
     memory[2346] = 32'd95;
     memory[2347] = 32'd168;
     memory[2348] = 32'd132;
     memory[2349] = 32'd212;
     memory[2350] = 32'd100;
     memory[2351] = 32'd146;
     memory[2352] = 32'd168;
     memory[2353] = 32'd183;
     memory[2354] = 32'd97;
     memory[2355] = 32'd164;
     memory[2356] = 32'd90;
     memory[2357] = 32'd137;
     memory[2358] = 32'd23;
     memory[2359] = 32'd87;
     memory[2360] = 32'd76;
     memory[2361] = 32'd231;
     memory[2362] = 32'd177;
     memory[2363] = 32'd244;
     memory[2364] = 32'd154;
     memory[2365] = 32'd215;
     memory[2366] = 32'd79;
     memory[2367] = 32'd230;
     memory[2368] = 32'd210;
     memory[2369] = 32'd123;
     memory[2370] = 32'd181;
     memory[2371] = 32'd23;
     memory[2372] = 32'd107;
     memory[2373] = 32'd91;
     memory[2374] = 32'd36;
     memory[2375] = 32'd221;
     memory[2376] = 32'd123;
     memory[2377] = 32'd105;
     memory[2378] = 32'd233;
     memory[2379] = 32'd231;
     memory[2380] = 32'd17;
     memory[2381] = 32'd81;
     memory[2382] = 32'd174;
     memory[2383] = 32'd84;
     memory[2384] = 32'd89;
     memory[2385] = 32'd212;
     memory[2386] = 32'd76;
     memory[2387] = 32'd205;
     memory[2388] = 32'd196;
     memory[2389] = 32'd162;
     memory[2390] = 32'd178;
     memory[2391] = 32'd32;
     memory[2392] = 32'd80;
     memory[2393] = 32'd207;
     memory[2394] = 32'd68;
     memory[2395] = 32'd11;
     memory[2396] = 32'd142;
     memory[2397] = 32'd82;
     memory[2398] = 32'd191;
     memory[2399] = 32'd139;
     memory[2400] = 32'd240;
     memory[2401] = 32'd15;
     memory[2402] = 32'd113;
     memory[2403] = 32'd6;
     memory[2404] = 32'd126;
     memory[2405] = 32'd10;
     memory[2406] = 32'd213;
     memory[2407] = 32'd192;
     memory[2408] = 32'd23;
     memory[2409] = 32'd118;
     memory[2410] = 32'd168;
     memory[2411] = 32'd198;
     memory[2412] = 32'd214;
     memory[2413] = 32'd20;
     memory[2414] = 32'd76;
     memory[2415] = 32'd163;
     memory[2416] = 32'd4;
     memory[2417] = 32'd51;
     memory[2418] = 32'd245;
     memory[2419] = 32'd123;
     memory[2420] = 32'd64;
     memory[2421] = 32'd183;
     memory[2422] = 32'd90;
     memory[2423] = 32'd48;
     memory[2424] = 32'd194;
     memory[2425] = 32'd154;
     memory[2426] = 32'd144;
     memory[2427] = 32'd128;
     memory[2428] = 32'd224;
     memory[2429] = 32'd90;
     memory[2430] = 32'd157;
     memory[2431] = 32'd174;
     memory[2432] = 32'd163;
     memory[2433] = 32'd209;
     memory[2434] = 32'd254;
     memory[2435] = 32'd65;
     memory[2436] = 32'd112;
     memory[2437] = 32'd21;
     memory[2438] = 32'd240;
     memory[2439] = 32'd18;
     memory[2440] = 32'd140;
     memory[2441] = 32'd129;
     memory[2442] = 32'd248;
     memory[2443] = 32'd71;
     memory[2444] = 32'd22;
     memory[2445] = 32'd219;
     memory[2446] = 32'd55;
     memory[2447] = 32'd25;
     memory[2448] = 32'd22;
     memory[2449] = 32'd168;
     memory[2450] = 32'd96;
     memory[2451] = 32'd97;
     memory[2452] = 32'd90;
     memory[2453] = 32'd117;
     memory[2454] = 32'd195;
     memory[2455] = 32'd198;
     memory[2456] = 32'd144;
     memory[2457] = 32'd77;
     memory[2458] = 32'd54;
     memory[2459] = 32'd200;
     memory[2460] = 32'd119;
     memory[2461] = 32'd19;
     memory[2462] = 32'd57;
     memory[2463] = 32'd104;
     memory[2464] = 32'd107;
     memory[2465] = 32'd222;
     memory[2466] = 32'd202;
     memory[2467] = 32'd47;
     memory[2468] = 32'd39;
     memory[2469] = 32'd217;
     memory[2470] = 32'd98;
     memory[2471] = 32'd247;
     memory[2472] = 32'd80;
     memory[2473] = 32'd237;
     memory[2474] = 32'd193;
     memory[2475] = 32'd87;
     memory[2476] = 32'd122;
     memory[2477] = 32'd87;
     memory[2478] = 32'd179;
     memory[2479] = 32'd99;
     memory[2480] = 32'd215;
     memory[2481] = 32'd40;
     memory[2482] = 32'd121;
     memory[2483] = 32'd181;
     memory[2484] = 32'd190;
     memory[2485] = 32'd69;
     memory[2486] = 32'd210;
     memory[2487] = 32'd4;
     memory[2488] = 32'd205;
     memory[2489] = 32'd124;
     memory[2490] = 32'd137;
     memory[2491] = 32'd116;
     memory[2492] = 32'd241;
     memory[2493] = 32'd145;
     memory[2494] = 32'd51;
     memory[2495] = 32'd213;
     memory[2496] = 32'd73;
     memory[2497] = 32'd145;
     memory[2498] = 32'd88;
     memory[2499] = 32'd44;
     memory[2500] = 32'd221;
     memory[2501] = 32'd127;
     memory[2502] = 32'd116;
     memory[2503] = 32'd201;
     memory[2504] = 32'd118;
     memory[2505] = 32'd125;
     memory[2506] = 32'd247;
     memory[2507] = 32'd222;
     memory[2508] = 32'd235;
     memory[2509] = 32'd7;
     memory[2510] = 32'd209;
     memory[2511] = 32'd44;
     memory[2512] = 32'd178;
     memory[2513] = 32'd159;
     memory[2514] = 32'd238;
     memory[2515] = 32'd26;
     memory[2516] = 32'd152;
     memory[2517] = 32'd216;
     memory[2518] = 32'd4;
     memory[2519] = 32'd158;
     memory[2520] = 32'd21;
     memory[2521] = 32'd82;
     memory[2522] = 32'd244;
     memory[2523] = 32'd39;
     memory[2524] = 32'd145;
     memory[2525] = 32'd69;
     memory[2526] = 32'd234;
     memory[2527] = 32'd5;
     memory[2528] = 32'd67;
     memory[2529] = 32'd119;
     memory[2530] = 32'd214;
     memory[2531] = 32'd201;
     memory[2532] = 32'd139;
     memory[2533] = 32'd254;
     memory[2534] = 32'd136;
     memory[2535] = 32'd182;
     memory[2536] = 32'd74;
     memory[2537] = 32'd213;
     memory[2538] = 32'd93;
     memory[2539] = 32'd11;
     memory[2540] = 32'd29;
     memory[2541] = 32'd90;
     memory[2542] = 32'd205;
     memory[2543] = 32'd178;
     memory[2544] = 32'd193;
     memory[2545] = 32'd67;
     memory[2546] = 32'd131;
     memory[2547] = 32'd4;
     memory[2548] = 32'd122;
     memory[2549] = 32'd3;
     memory[2550] = 32'd156;
     memory[2551] = 32'd168;
     memory[2552] = 32'd50;
     memory[2553] = 32'd211;
     memory[2554] = 32'd163;
     memory[2555] = 32'd97;
     memory[2556] = 32'd180;
     memory[2557] = 32'd73;
     memory[2558] = 32'd30;
     memory[2559] = 32'd229;
     memory[2560] = 32'd139;
     memory[2561] = 32'd97;
     memory[2562] = 32'd20;
     memory[2563] = 32'd93;
     memory[2564] = 32'd198;
     memory[2565] = 32'd116;
     memory[2566] = 32'd24;
     memory[2567] = 32'd171;
     memory[2568] = 32'd6;
     memory[2569] = 32'd74;
     memory[2570] = 32'd173;
     memory[2571] = 32'd6;
     memory[2572] = 32'd64;
     memory[2573] = 32'd211;
     memory[2574] = 32'd228;
     memory[2575] = 32'd240;
     memory[2576] = 32'd88;
     memory[2577] = 32'd44;
     memory[2578] = 32'd124;
     memory[2579] = 32'd99;
     memory[2580] = 32'd4;
     memory[2581] = 32'd218;
     memory[2582] = 32'd104;
     memory[2583] = 32'd203;
     memory[2584] = 32'd115;
     memory[2585] = 32'd35;
     memory[2586] = 32'd148;
     memory[2587] = 32'd14;
     memory[2588] = 32'd154;
     memory[2589] = 32'd23;
     memory[2590] = 32'd4;
     memory[2591] = 32'd115;
     memory[2592] = 32'd158;
     memory[2593] = 32'd158;
     memory[2594] = 32'd231;
     memory[2595] = 32'd6;
     memory[2596] = 32'd150;
     memory[2597] = 32'd123;
     memory[2598] = 32'd167;
     memory[2599] = 32'd212;
     memory[2600] = 32'd9;
     memory[2601] = 32'd129;
     memory[2602] = 32'd96;
     memory[2603] = 32'd134;
     memory[2604] = 32'd6;
     memory[2605] = 32'd245;
     memory[2606] = 32'd250;
     memory[2607] = 32'd145;
     memory[2608] = 32'd2;
     memory[2609] = 32'd75;
     memory[2610] = 32'd123;
     memory[2611] = 32'd148;
     memory[2612] = 32'd141;
     memory[2613] = 32'd240;
     memory[2614] = 32'd128;
     memory[2615] = 32'd235;
     memory[2616] = 32'd229;
     memory[2617] = 32'd15;
     memory[2618] = 32'd41;
     memory[2619] = 32'd121;
     memory[2620] = 32'd34;
     memory[2621] = 32'd166;
     memory[2622] = 32'd214;
     memory[2623] = 32'd26;
     memory[2624] = 32'd158;
     memory[2625] = 32'd245;
     memory[2626] = 32'd237;
     memory[2627] = 32'd249;
     memory[2628] = 32'd173;
     memory[2629] = 32'd224;
     memory[2630] = 32'd58;
     memory[2631] = 32'd236;
     memory[2632] = 32'd8;
     memory[2633] = 32'd244;
     memory[2634] = 32'd122;
     memory[2635] = 32'd74;
     memory[2636] = 32'd131;
     memory[2637] = 32'd188;
     memory[2638] = 32'd67;
     memory[2639] = 32'd149;
     memory[2640] = 32'd136;
     memory[2641] = 32'd245;
     memory[2642] = 32'd42;
     memory[2643] = 32'd224;
     memory[2644] = 32'd126;
     memory[2645] = 32'd76;
     memory[2646] = 32'd80;
     memory[2647] = 32'd105;
     memory[2648] = 32'd97;
     memory[2649] = 32'd145;
     memory[2650] = 32'd208;
     memory[2651] = 32'd88;
     memory[2652] = 32'd230;
     memory[2653] = 32'd126;
     memory[2654] = 32'd246;
     memory[2655] = 32'd237;
     memory[2656] = 32'd152;
     memory[2657] = 32'd24;
     memory[2658] = 32'd218;
     memory[2659] = 32'd39;
     memory[2660] = 32'd84;
     memory[2661] = 32'd107;
     memory[2662] = 32'd36;
     memory[2663] = 32'd55;
     memory[2664] = 32'd118;
     memory[2665] = 32'd160;
     memory[2666] = 32'd173;
     memory[2667] = 32'd182;
     memory[2668] = 32'd53;
     memory[2669] = 32'd146;
     memory[2670] = 32'd131;
     memory[2671] = 32'd164;
     memory[2672] = 32'd58;
     memory[2673] = 32'd14;
     memory[2674] = 32'd76;
     memory[2675] = 32'd136;
     memory[2676] = 32'd110;
     memory[2677] = 32'd68;
     memory[2678] = 32'd207;
     memory[2679] = 32'd181;
     memory[2680] = 32'd171;
     memory[2681] = 32'd142;
     memory[2682] = 32'd237;
     memory[2683] = 32'd129;
     memory[2684] = 32'd204;
     memory[2685] = 32'd227;
     memory[2686] = 32'd16;
     memory[2687] = 32'd5;
     memory[2688] = 32'd92;
     memory[2689] = 32'd145;
     memory[2690] = 32'd3;
     memory[2691] = 32'd9;
     memory[2692] = 32'd19;
     memory[2693] = 32'd106;
     memory[2694] = 32'd90;
     memory[2695] = 32'd8;
     memory[2696] = 32'd98;
     memory[2697] = 32'd75;
     memory[2698] = 32'd6;
     memory[2699] = 32'd220;
     memory[2700] = 32'd139;
     memory[2701] = 32'd106;
     memory[2702] = 32'd165;
     memory[2703] = 32'd243;
     memory[2704] = 32'd131;
     memory[2705] = 32'd225;
     memory[2706] = 32'd59;
     memory[2707] = 32'd103;
     memory[2708] = 32'd56;
     memory[2709] = 32'd185;
     memory[2710] = 32'd159;
     memory[2711] = 32'd71;
     memory[2712] = 32'd156;
     memory[2713] = 32'd42;
     memory[2714] = 32'd75;
     memory[2715] = 32'd60;
     memory[2716] = 32'd167;
     memory[2717] = 32'd249;
     memory[2718] = 32'd120;
     memory[2719] = 32'd55;
     memory[2720] = 32'd190;
     memory[2721] = 32'd164;
     memory[2722] = 32'd96;
     memory[2723] = 32'd72;
     memory[2724] = 32'd123;
     memory[2725] = 32'd123;
     memory[2726] = 32'd32;
     memory[2727] = 32'd6;
     memory[2728] = 32'd190;
     memory[2729] = 32'd155;
     memory[2730] = 32'd48;
     memory[2731] = 32'd214;
     memory[2732] = 32'd207;
     memory[2733] = 32'd171;
     memory[2734] = 32'd149;
     memory[2735] = 32'd219;
     memory[2736] = 32'd96;
     memory[2737] = 32'd234;
     memory[2738] = 32'd253;
     memory[2739] = 32'd178;
     memory[2740] = 32'd190;
     memory[2741] = 32'd230;
     memory[2742] = 32'd10;
     memory[2743] = 32'd207;
     memory[2744] = 32'd29;
     memory[2745] = 32'd208;
     memory[2746] = 32'd246;
     memory[2747] = 32'd220;
     memory[2748] = 32'd219;
     memory[2749] = 32'd217;
     memory[2750] = 32'd85;
     memory[2751] = 32'd19;
     memory[2752] = 32'd163;
     memory[2753] = 32'd236;
     memory[2754] = 32'd87;
     memory[2755] = 32'd22;
     memory[2756] = 32'd92;
     memory[2757] = 32'd249;
     memory[2758] = 32'd4;
     memory[2759] = 32'd103;
     memory[2760] = 32'd105;
     memory[2761] = 32'd16;
     memory[2762] = 32'd131;
     memory[2763] = 32'd118;
     memory[2764] = 32'd206;
     memory[2765] = 32'd126;
     memory[2766] = 32'd103;
     memory[2767] = 32'd179;
     memory[2768] = 32'd254;
     memory[2769] = 32'd0;
     memory[2770] = 32'd81;
     memory[2771] = 32'd181;
     memory[2772] = 32'd85;
     memory[2773] = 32'd84;
     memory[2774] = 32'd37;
     memory[2775] = 32'd148;
     memory[2776] = 32'd51;
     memory[2777] = 32'd144;
     memory[2778] = 32'd215;
     memory[2779] = 32'd237;
     memory[2780] = 32'd68;
     memory[2781] = 32'd49;
     memory[2782] = 32'd58;
     memory[2783] = 32'd179;
     memory[2784] = 32'd140;
     memory[2785] = 32'd229;
     memory[2786] = 32'd89;
     memory[2787] = 32'd224;
     memory[2788] = 32'd7;
     memory[2789] = 32'd89;
     memory[2790] = 32'd176;
     memory[2791] = 32'd38;
     memory[2792] = 32'd229;
     memory[2793] = 32'd4;
     memory[2794] = 32'd157;
     memory[2795] = 32'd32;
     memory[2796] = 32'd57;
     memory[2797] = 32'd246;
     memory[2798] = 32'd127;
     memory[2799] = 32'd210;
     memory[2800] = 32'd86;
     memory[2801] = 32'd208;
     memory[2802] = 32'd93;
     memory[2803] = 32'd114;
     memory[2804] = 32'd252;
     memory[2805] = 32'd54;
     memory[2806] = 32'd101;
     memory[2807] = 32'd90;
     memory[2808] = 32'd222;
     memory[2809] = 32'd239;
     memory[2810] = 32'd225;
     memory[2811] = 32'd14;
     memory[2812] = 32'd227;
     memory[2813] = 32'd123;
     memory[2814] = 32'd40;
     memory[2815] = 32'd219;
     memory[2816] = 32'd148;
     memory[2817] = 32'd253;
     memory[2818] = 32'd190;
     memory[2819] = 32'd85;
     memory[2820] = 32'd31;
     memory[2821] = 32'd116;
     memory[2822] = 32'd153;
     memory[2823] = 32'd120;
     memory[2824] = 32'd34;
     memory[2825] = 32'd51;
     memory[2826] = 32'd247;
     memory[2827] = 32'd169;
     memory[2828] = 32'd203;
     memory[2829] = 32'd163;
     memory[2830] = 32'd191;
     memory[2831] = 32'd153;
     memory[2832] = 32'd248;
     memory[2833] = 32'd226;
     memory[2834] = 32'd78;
     memory[2835] = 32'd120;
     memory[2836] = 32'd46;
     memory[2837] = 32'd146;
     memory[2838] = 32'd89;
     memory[2839] = 32'd90;
     memory[2840] = 32'd225;
     memory[2841] = 32'd147;
     memory[2842] = 32'd252;
     memory[2843] = 32'd30;
     memory[2844] = 32'd149;
     memory[2845] = 32'd134;
     memory[2846] = 32'd38;
     memory[2847] = 32'd80;
     memory[2848] = 32'd73;
     memory[2849] = 32'd41;
     memory[2850] = 32'd185;
     memory[2851] = 32'd169;
     memory[2852] = 32'd35;
     memory[2853] = 32'd178;
     memory[2854] = 32'd62;
     memory[2855] = 32'd249;
     memory[2856] = 32'd66;
     memory[2857] = 32'd182;
     memory[2858] = 32'd99;
     memory[2859] = 32'd149;
     memory[2860] = 32'd145;
     memory[2861] = 32'd27;
     memory[2862] = 32'd219;
     memory[2863] = 32'd186;
     memory[2864] = 32'd104;
     memory[2865] = 32'd231;
     memory[2866] = 32'd202;
     memory[2867] = 32'd71;
     memory[2868] = 32'd131;
     memory[2869] = 32'd4;
     memory[2870] = 32'd88;
     memory[2871] = 32'd25;
     memory[2872] = 32'd188;
     memory[2873] = 32'd0;
     memory[2874] = 32'd156;
     memory[2875] = 32'd235;
     memory[2876] = 32'd32;
     memory[2877] = 32'd224;
     memory[2878] = 32'd21;
     memory[2879] = 32'd112;
     memory[2880] = 32'd69;
     memory[2881] = 32'd86;
     memory[2882] = 32'd121;
     memory[2883] = 32'd226;
     memory[2884] = 32'd221;
     memory[2885] = 32'd117;
     memory[2886] = 32'd242;
     memory[2887] = 32'd12;
     memory[2888] = 32'd202;
     memory[2889] = 32'd190;
     memory[2890] = 32'd211;
     memory[2891] = 32'd209;
     memory[2892] = 32'd79;
     memory[2893] = 32'd124;
     memory[2894] = 32'd32;
     memory[2895] = 32'd224;
     memory[2896] = 32'd7;
     memory[2897] = 32'd5;
     memory[2898] = 32'd204;
     memory[2899] = 32'd6;
     memory[2900] = 32'd136;
     memory[2901] = 32'd253;
     memory[2902] = 32'd53;
     memory[2903] = 32'd4;
     memory[2904] = 32'd58;
     memory[2905] = 32'd72;
     memory[2906] = 32'd51;
     memory[2907] = 32'd32;
     memory[2908] = 32'd219;
     memory[2909] = 32'd197;
     memory[2910] = 32'd187;
     memory[2911] = 32'd221;
     memory[2912] = 32'd14;
     memory[2913] = 32'd14;
     memory[2914] = 32'd242;
     memory[2915] = 32'd189;
     memory[2916] = 32'd180;
     memory[2917] = 32'd228;
     memory[2918] = 32'd41;
     memory[2919] = 32'd136;
     memory[2920] = 32'd172;
     memory[2921] = 32'd37;
     memory[2922] = 32'd64;
     memory[2923] = 32'd116;
     memory[2924] = 32'd224;
     memory[2925] = 32'd11;
     memory[2926] = 32'd103;
     memory[2927] = 32'd226;
     memory[2928] = 32'd178;
     memory[2929] = 32'd94;
     memory[2930] = 32'd87;
     memory[2931] = 32'd55;
     memory[2932] = 32'd110;
     memory[2933] = 32'd147;
     memory[2934] = 32'd122;
     memory[2935] = 32'd53;
     memory[2936] = 32'd180;
     memory[2937] = 32'd92;
     memory[2938] = 32'd18;
     memory[2939] = 32'd227;
     memory[2940] = 32'd2;
     memory[2941] = 32'd169;
     memory[2942] = 32'd207;
     memory[2943] = 32'd205;
     memory[2944] = 32'd43;
     memory[2945] = 32'd140;
     memory[2946] = 32'd120;
     memory[2947] = 32'd167;
     memory[2948] = 32'd39;
     memory[2949] = 32'd183;
     memory[2950] = 32'd229;
     memory[2951] = 32'd110;
     memory[2952] = 32'd245;
     memory[2953] = 32'd122;
     memory[2954] = 32'd41;
     memory[2955] = 32'd152;
     memory[2956] = 32'd241;
     memory[2957] = 32'd202;
     memory[2958] = 32'd215;
     memory[2959] = 32'd66;
     memory[2960] = 32'd79;
     memory[2961] = 32'd93;
     memory[2962] = 32'd106;
     memory[2963] = 32'd29;
     memory[2964] = 32'd120;
     memory[2965] = 32'd208;
     memory[2966] = 32'd83;
     memory[2967] = 32'd1;
     memory[2968] = 32'd89;
     memory[2969] = 32'd136;
     memory[2970] = 32'd82;
     memory[2971] = 32'd222;
     memory[2972] = 32'd124;
     memory[2973] = 32'd20;
     memory[2974] = 32'd106;
     memory[2975] = 32'd38;
     memory[2976] = 32'd147;
     memory[2977] = 32'd149;
     memory[2978] = 32'd120;
     memory[2979] = 32'd162;
     memory[2980] = 32'd93;
     memory[2981] = 32'd32;
     memory[2982] = 32'd132;
     memory[2983] = 32'd212;
     memory[2984] = 32'd199;
     memory[2985] = 32'd20;
     memory[2986] = 32'd236;
     memory[2987] = 32'd119;
     memory[2988] = 32'd9;
     memory[2989] = 32'd155;
     memory[2990] = 32'd101;
     memory[2991] = 32'd100;
     memory[2992] = 32'd155;
     memory[2993] = 32'd96;
     memory[2994] = 32'd63;
     memory[2995] = 32'd171;
     memory[2996] = 32'd242;
     memory[2997] = 32'd186;
     memory[2998] = 32'd216;
     memory[2999] = 32'd230;
     memory[3000] = 32'd70;
     memory[3001] = 32'd159;
     memory[3002] = 32'd59;
     memory[3003] = 32'd222;
     memory[3004] = 32'd22;
     memory[3005] = 32'd155;
     memory[3006] = 32'd223;
     memory[3007] = 32'd125;
     memory[3008] = 32'd25;
     memory[3009] = 32'd23;
     memory[3010] = 32'd107;
     memory[3011] = 32'd84;
     memory[3012] = 32'd70;
     memory[3013] = 32'd110;
     memory[3014] = 32'd2;
     memory[3015] = 32'd225;
     memory[3016] = 32'd171;
     memory[3017] = 32'd58;
     memory[3018] = 32'd22;
     memory[3019] = 32'd72;
     memory[3020] = 32'd181;
     memory[3021] = 32'd21;
     memory[3022] = 32'd134;
     memory[3023] = 32'd232;
     memory[3024] = 32'd68;
     memory[3025] = 32'd70;
     memory[3026] = 32'd13;
     memory[3027] = 32'd55;
     memory[3028] = 32'd107;
     memory[3029] = 32'd64;
     memory[3030] = 32'd243;
     memory[3031] = 32'd76;
     memory[3032] = 32'd105;
     memory[3033] = 32'd60;
     memory[3034] = 32'd241;
     memory[3035] = 32'd204;
     memory[3036] = 32'd31;
     memory[3037] = 32'd0;
     memory[3038] = 32'd14;
     memory[3039] = 32'd243;
     memory[3040] = 32'd161;
     memory[3041] = 32'd26;
     memory[3042] = 32'd243;
     memory[3043] = 32'd232;
     memory[3044] = 32'd38;
     memory[3045] = 32'd219;
     memory[3046] = 32'd55;
     memory[3047] = 32'd30;
     memory[3048] = 32'd171;
     memory[3049] = 32'd144;
     memory[3050] = 32'd168;
     memory[3051] = 32'd178;
     memory[3052] = 32'd62;
     memory[3053] = 32'd191;
     memory[3054] = 32'd26;
     memory[3055] = 32'd117;
     memory[3056] = 32'd183;
     memory[3057] = 32'd30;
     memory[3058] = 32'd197;
     memory[3059] = 32'd51;
     memory[3060] = 32'd234;
     memory[3061] = 32'd93;
     memory[3062] = 32'd240;
     memory[3063] = 32'd253;
     memory[3064] = 32'd113;
     memory[3065] = 32'd24;
     memory[3066] = 32'd83;
     memory[3067] = 32'd130;
     memory[3068] = 32'd153;
     memory[3069] = 32'd46;
     memory[3070] = 32'd30;
     memory[3071] = 32'd235;
     memory[3072] = 32'd212;
     memory[3073] = 32'd218;
     memory[3074] = 32'd33;
     memory[3075] = 32'd150;
     memory[3076] = 32'd53;
     memory[3077] = 32'd33;
     memory[3078] = 32'd49;
     memory[3079] = 32'd229;
     memory[3080] = 32'd38;
     memory[3081] = 32'd124;
     memory[3082] = 32'd159;
     memory[3083] = 32'd86;
     memory[3084] = 32'd222;
     memory[3085] = 32'd136;
     memory[3086] = 32'd10;
     memory[3087] = 32'd150;
     memory[3088] = 32'd161;
     memory[3089] = 32'd85;
     memory[3090] = 32'd216;
     memory[3091] = 32'd141;
     memory[3092] = 32'd124;
     memory[3093] = 32'd134;
     memory[3094] = 32'd184;
     memory[3095] = 32'd41;
     memory[3096] = 32'd67;
     memory[3097] = 32'd45;
     memory[3098] = 32'd87;
     memory[3099] = 32'd156;
     memory[3100] = 32'd170;
     memory[3101] = 32'd147;
     memory[3102] = 32'd78;
     memory[3103] = 32'd41;
     memory[3104] = 32'd208;
     memory[3105] = 32'd102;
     memory[3106] = 32'd226;
     memory[3107] = 32'd97;
     memory[3108] = 32'd208;
     memory[3109] = 32'd202;
     memory[3110] = 32'd59;
     memory[3111] = 32'd46;
     memory[3112] = 32'd106;
     memory[3113] = 32'd198;
     memory[3114] = 32'd6;
     memory[3115] = 32'd23;
     memory[3116] = 32'd223;
     memory[3117] = 32'd73;
     memory[3118] = 32'd177;
     memory[3119] = 32'd251;
     memory[3120] = 32'd140;
     memory[3121] = 32'd61;
     memory[3122] = 32'd239;
     memory[3123] = 32'd250;
     memory[3124] = 32'd85;
     memory[3125] = 32'd214;
     memory[3126] = 32'd213;
     memory[3127] = 32'd247;
     memory[3128] = 32'd68;
     memory[3129] = 32'd121;
     memory[3130] = 32'd191;
     memory[3131] = 32'd14;
     memory[3132] = 32'd38;
     memory[3133] = 32'd121;
     memory[3134] = 32'd0;
     memory[3135] = 32'd113;
     memory[3136] = 32'd16;
     memory[3137] = 32'd46;
     memory[3138] = 32'd153;
     memory[3139] = 32'd75;
     memory[3140] = 32'd247;
     memory[3141] = 32'd103;
     memory[3142] = 32'd201;
     memory[3143] = 32'd45;
     memory[3144] = 32'd102;
     memory[3145] = 32'd121;
     memory[3146] = 32'd144;
     memory[3147] = 32'd97;
     memory[3148] = 32'd153;
     memory[3149] = 32'd2;
     memory[3150] = 32'd87;
     memory[3151] = 32'd204;
     memory[3152] = 32'd168;
     memory[3153] = 32'd54;
     memory[3154] = 32'd24;
     memory[3155] = 32'd185;
     memory[3156] = 32'd54;
     memory[3157] = 32'd80;
     memory[3158] = 32'd238;
     memory[3159] = 32'd159;
     memory[3160] = 32'd141;
     memory[3161] = 32'd49;
     memory[3162] = 32'd181;
     memory[3163] = 32'd187;
     memory[3164] = 32'd103;
     memory[3165] = 32'd209;
     memory[3166] = 32'd183;
     memory[3167] = 32'd155;
     memory[3168] = 32'd131;
     memory[3169] = 32'd248;
     memory[3170] = 32'd253;
     memory[3171] = 32'd158;
     memory[3172] = 32'd122;
     memory[3173] = 32'd117;
     memory[3174] = 32'd229;
     memory[3175] = 32'd212;
     memory[3176] = 32'd66;
     memory[3177] = 32'd48;
     memory[3178] = 32'd29;
     memory[3179] = 32'd210;
     memory[3180] = 32'd217;
     memory[3181] = 32'd62;
     memory[3182] = 32'd72;
     memory[3183] = 32'd21;
     memory[3184] = 32'd187;
     memory[3185] = 32'd137;
     memory[3186] = 32'd253;
     memory[3187] = 32'd133;
     memory[3188] = 32'd156;
     memory[3189] = 32'd156;
     memory[3190] = 32'd144;
     memory[3191] = 32'd93;
     memory[3192] = 32'd206;
     memory[3193] = 32'd212;
     memory[3194] = 32'd180;
     memory[3195] = 32'd197;
     memory[3196] = 32'd36;
     memory[3197] = 32'd208;
     memory[3198] = 32'd231;
     memory[3199] = 32'd4;
     memory[3200] = 32'd110;
     memory[3201] = 32'd198;
     memory[3202] = 32'd96;
     memory[3203] = 32'd244;
     memory[3204] = 32'd5;
     memory[3205] = 32'd14;
     memory[3206] = 32'd0;
     memory[3207] = 32'd163;
     memory[3208] = 32'd63;
     memory[3209] = 32'd253;
     memory[3210] = 32'd184;
     memory[3211] = 32'd65;
     memory[3212] = 32'd189;
     memory[3213] = 32'd61;
     memory[3214] = 32'd2;
     memory[3215] = 32'd104;
     memory[3216] = 32'd254;
     memory[3217] = 32'd157;
     memory[3218] = 32'd108;
     memory[3219] = 32'd211;
     memory[3220] = 32'd175;
     memory[3221] = 32'd28;
     memory[3222] = 32'd54;
     memory[3223] = 32'd66;
     memory[3224] = 32'd235;
     memory[3225] = 32'd172;
     memory[3226] = 32'd23;
     memory[3227] = 32'd107;
     memory[3228] = 32'd87;
     memory[3229] = 32'd31;
     memory[3230] = 32'd196;
     memory[3231] = 32'd42;
     memory[3232] = 32'd223;
     memory[3233] = 32'd78;
     memory[3234] = 32'd121;
     memory[3235] = 32'd196;
     memory[3236] = 32'd70;
     memory[3237] = 32'd252;
     memory[3238] = 32'd68;
     memory[3239] = 32'd223;
     memory[3240] = 32'd179;
     memory[3241] = 32'd215;
     memory[3242] = 32'd18;
     memory[3243] = 32'd92;
     memory[3244] = 32'd5;
     memory[3245] = 32'd107;
     memory[3246] = 32'd65;
     memory[3247] = 32'd137;
     memory[3248] = 32'd69;
     memory[3249] = 32'd94;
     memory[3250] = 32'd51;
     memory[3251] = 32'd235;
     memory[3252] = 32'd173;
     memory[3253] = 32'd100;
     memory[3254] = 32'd221;
     memory[3255] = 32'd208;
     memory[3256] = 32'd183;
     memory[3257] = 32'd108;
     memory[3258] = 32'd157;
     memory[3259] = 32'd210;
     memory[3260] = 32'd169;
     memory[3261] = 32'd218;
     memory[3262] = 32'd42;
     memory[3263] = 32'd62;
     memory[3264] = 32'd27;
     memory[3265] = 32'd241;
     memory[3266] = 32'd211;
     memory[3267] = 32'd155;
     memory[3268] = 32'd242;
     memory[3269] = 32'd126;
     memory[3270] = 32'd209;
     memory[3271] = 32'd92;
     memory[3272] = 32'd66;
     memory[3273] = 32'd51;
     memory[3274] = 32'd132;
     memory[3275] = 32'd217;
     memory[3276] = 32'd202;
     memory[3277] = 32'd187;
     memory[3278] = 32'd68;
     memory[3279] = 32'd11;
     memory[3280] = 32'd33;
     memory[3281] = 32'd130;
     memory[3282] = 32'd172;
     memory[3283] = 32'd17;
     memory[3284] = 32'd247;
     memory[3285] = 32'd18;
     memory[3286] = 32'd188;
     memory[3287] = 32'd161;
     memory[3288] = 32'd192;
     memory[3289] = 32'd208;
     memory[3290] = 32'd45;
     memory[3291] = 32'd164;
     memory[3292] = 32'd234;
     memory[3293] = 32'd178;
     memory[3294] = 32'd156;
     memory[3295] = 32'd195;
     memory[3296] = 32'd133;
     memory[3297] = 32'd50;
     memory[3298] = 32'd26;
     memory[3299] = 32'd242;
     memory[3300] = 32'd54;
     memory[3301] = 32'd102;
     memory[3302] = 32'd147;
     memory[3303] = 32'd184;
     memory[3304] = 32'd6;
     memory[3305] = 32'd230;
     memory[3306] = 32'd122;
     memory[3307] = 32'd204;
     memory[3308] = 32'd28;
     memory[3309] = 32'd2;
     memory[3310] = 32'd0;
     memory[3311] = 32'd16;
     memory[3312] = 32'd51;
     memory[3313] = 32'd222;
     memory[3314] = 32'd244;
     memory[3315] = 32'd120;
     memory[3316] = 32'd148;
     memory[3317] = 32'd24;
     memory[3318] = 32'd8;
     memory[3319] = 32'd39;
     memory[3320] = 32'd249;
     memory[3321] = 32'd171;
     memory[3322] = 32'd245;
     memory[3323] = 32'd193;
     memory[3324] = 32'd234;
     memory[3325] = 32'd178;
     memory[3326] = 32'd0;
     memory[3327] = 32'd128;
     memory[3328] = 32'd193;
     memory[3329] = 32'd240;
     memory[3330] = 32'd16;
     memory[3331] = 32'd254;
     memory[3332] = 32'd79;
     memory[3333] = 32'd197;
     memory[3334] = 32'd131;
     memory[3335] = 32'd95;
     memory[3336] = 32'd195;
     memory[3337] = 32'd250;
     memory[3338] = 32'd21;
     memory[3339] = 32'd9;
     memory[3340] = 32'd187;
     memory[3341] = 32'd216;
     memory[3342] = 32'd108;
     memory[3343] = 32'd237;
     memory[3344] = 32'd16;
     memory[3345] = 32'd232;
     memory[3346] = 32'd77;
     memory[3347] = 32'd23;
     memory[3348] = 32'd216;
     memory[3349] = 32'd33;
     memory[3350] = 32'd62;
     memory[3351] = 32'd233;
     memory[3352] = 32'd251;
     memory[3353] = 32'd113;
     memory[3354] = 32'd198;
     memory[3355] = 32'd50;
     memory[3356] = 32'd101;
     memory[3357] = 32'd111;
     memory[3358] = 32'd69;
     memory[3359] = 32'd54;
     memory[3360] = 32'd230;
     memory[3361] = 32'd23;
     memory[3362] = 32'd185;
     memory[3363] = 32'd214;
     memory[3364] = 32'd173;
     memory[3365] = 32'd143;
     memory[3366] = 32'd205;
     memory[3367] = 32'd172;
     memory[3368] = 32'd40;
     memory[3369] = 32'd179;
     memory[3370] = 32'd241;
     memory[3371] = 32'd30;
     memory[3372] = 32'd224;
     memory[3373] = 32'd228;
     memory[3374] = 32'd234;
     memory[3375] = 32'd154;
     memory[3376] = 32'd158;
     memory[3377] = 32'd167;
     memory[3378] = 32'd216;
     memory[3379] = 32'd184;
     memory[3380] = 32'd147;
     memory[3381] = 32'd64;
     memory[3382] = 32'd165;
     memory[3383] = 32'd203;
     memory[3384] = 32'd103;
     memory[3385] = 32'd156;
     memory[3386] = 32'd173;
     memory[3387] = 32'd96;
     memory[3388] = 32'd214;
     memory[3389] = 32'd153;
     memory[3390] = 32'd180;
     memory[3391] = 32'd207;
     memory[3392] = 32'd80;
     memory[3393] = 32'd228;
     memory[3394] = 32'd98;
     memory[3395] = 32'd88;
     memory[3396] = 32'd0;
     memory[3397] = 32'd144;
     memory[3398] = 32'd12;
     memory[3399] = 32'd190;
     memory[3400] = 32'd45;
     memory[3401] = 32'd102;
     memory[3402] = 32'd205;
     memory[3403] = 32'd188;
     memory[3404] = 32'd22;
     memory[3405] = 32'd233;
     memory[3406] = 32'd55;
     memory[3407] = 32'd201;
     memory[3408] = 32'd209;
     memory[3409] = 32'd139;
     memory[3410] = 32'd230;
     memory[3411] = 32'd135;
     memory[3412] = 32'd97;
     memory[3413] = 32'd228;
     memory[3414] = 32'd206;
     memory[3415] = 32'd20;
     memory[3416] = 32'd40;
     memory[3417] = 32'd193;
     memory[3418] = 32'd233;
     memory[3419] = 32'd152;
     memory[3420] = 32'd132;
     memory[3421] = 32'd44;
     memory[3422] = 32'd168;
     memory[3423] = 32'd216;
     memory[3424] = 32'd177;
     memory[3425] = 32'd138;
     memory[3426] = 32'd6;
     memory[3427] = 32'd222;
     memory[3428] = 32'd142;
     memory[3429] = 32'd67;
     memory[3430] = 32'd213;
     memory[3431] = 32'd49;
     memory[3432] = 32'd150;
     memory[3433] = 32'd147;
     memory[3434] = 32'd224;
     memory[3435] = 32'd64;
     memory[3436] = 32'd165;
     memory[3437] = 32'd119;
     memory[3438] = 32'd240;
     memory[3439] = 32'd84;
     memory[3440] = 32'd82;
     memory[3441] = 32'd135;
     memory[3442] = 32'd42;
     memory[3443] = 32'd188;
     memory[3444] = 32'd44;
     memory[3445] = 32'd60;
     memory[3446] = 32'd198;
     memory[3447] = 32'd190;
     memory[3448] = 32'd76;
     memory[3449] = 32'd121;
     memory[3450] = 32'd170;
     memory[3451] = 32'd210;
     memory[3452] = 32'd213;
     memory[3453] = 32'd105;
     memory[3454] = 32'd101;
     memory[3455] = 32'd71;
     memory[3456] = 32'd198;
     memory[3457] = 32'd94;
     memory[3458] = 32'd243;
     memory[3459] = 32'd193;
     memory[3460] = 32'd221;
     memory[3461] = 32'd215;
     memory[3462] = 32'd144;
     memory[3463] = 32'd101;
     memory[3464] = 32'd9;
     memory[3465] = 32'd189;
     memory[3466] = 32'd154;
     memory[3467] = 32'd237;
     memory[3468] = 32'd106;
     memory[3469] = 32'd174;
     memory[3470] = 32'd55;
     memory[3471] = 32'd162;
     memory[3472] = 32'd69;
     memory[3473] = 32'd84;
     memory[3474] = 32'd167;
     memory[3475] = 32'd114;
     memory[3476] = 32'd123;
     memory[3477] = 32'd162;
     memory[3478] = 32'd8;
     memory[3479] = 32'd7;
     memory[3480] = 32'd8;
     memory[3481] = 32'd134;
     memory[3482] = 32'd252;
     memory[3483] = 32'd55;
     memory[3484] = 32'd250;
     memory[3485] = 32'd108;
     memory[3486] = 32'd41;
     memory[3487] = 32'd202;
     memory[3488] = 32'd89;
     memory[3489] = 32'd239;
     memory[3490] = 32'd71;
     memory[3491] = 32'd181;
     memory[3492] = 32'd108;
     memory[3493] = 32'd166;
     memory[3494] = 32'd141;
     memory[3495] = 32'd88;
     memory[3496] = 32'd34;
     memory[3497] = 32'd157;
     memory[3498] = 32'd234;
     memory[3499] = 32'd28;
     memory[3500] = 32'd99;
     memory[3501] = 32'd63;
     memory[3502] = 32'd97;
     memory[3503] = 32'd13;
     memory[3504] = 32'd224;
     memory[3505] = 32'd176;
     memory[3506] = 32'd147;
     memory[3507] = 32'd35;
     memory[3508] = 32'd237;
     memory[3509] = 32'd251;
     memory[3510] = 32'd138;
     memory[3511] = 32'd137;
     memory[3512] = 32'd8;
     memory[3513] = 32'd97;
     memory[3514] = 32'd252;
     memory[3515] = 32'd134;
     memory[3516] = 32'd140;
     memory[3517] = 32'd71;
     memory[3518] = 32'd162;
     memory[3519] = 32'd199;
     memory[3520] = 32'd220;
     memory[3521] = 32'd244;
     memory[3522] = 32'd46;
     memory[3523] = 32'd150;
     memory[3524] = 32'd106;
     memory[3525] = 32'd244;
     memory[3526] = 32'd201;
     memory[3527] = 32'd218;
     memory[3528] = 32'd56;
     memory[3529] = 32'd21;
     memory[3530] = 32'd158;
     memory[3531] = 32'd101;
     memory[3532] = 32'd169;
     memory[3533] = 32'd249;
     memory[3534] = 32'd148;
     memory[3535] = 32'd132;
     memory[3536] = 32'd56;
     memory[3537] = 32'd186;
     memory[3538] = 32'd219;
     memory[3539] = 32'd172;
     memory[3540] = 32'd114;
     memory[3541] = 32'd92;
     memory[3542] = 32'd111;
     memory[3543] = 32'd52;
     memory[3544] = 32'd211;
     memory[3545] = 32'd169;
     memory[3546] = 32'd247;
     memory[3547] = 32'd237;
     memory[3548] = 32'd9;
     memory[3549] = 32'd151;
     memory[3550] = 32'd161;
     memory[3551] = 32'd52;
     memory[3552] = 32'd161;
     memory[3553] = 32'd204;
     memory[3554] = 32'd221;
     memory[3555] = 32'd127;
     memory[3556] = 32'd166;
     memory[3557] = 32'd195;
     memory[3558] = 32'd115;
     memory[3559] = 32'd193;
     memory[3560] = 32'd63;
     memory[3561] = 32'd137;
     memory[3562] = 32'd175;
     memory[3563] = 32'd210;
     memory[3564] = 32'd2;
     memory[3565] = 32'd54;
     memory[3566] = 32'd71;
     memory[3567] = 32'd216;
     memory[3568] = 32'd138;
     memory[3569] = 32'd232;
     memory[3570] = 32'd201;
     memory[3571] = 32'd202;
     memory[3572] = 32'd184;
     memory[3573] = 32'd144;
     memory[3574] = 32'd231;
     memory[3575] = 32'd139;
     memory[3576] = 32'd73;
     memory[3577] = 32'd17;
     memory[3578] = 32'd190;
     memory[3579] = 32'd236;
     memory[3580] = 32'd153;
     memory[3581] = 32'd214;
     memory[3582] = 32'd140;
     memory[3583] = 32'd66;
     memory[3584] = 32'd72;
     memory[3585] = 32'd148;
     memory[3586] = 32'd170;
     memory[3587] = 32'd144;
     memory[3588] = 32'd25;
     memory[3589] = 32'd138;
     memory[3590] = 32'd76;
     memory[3591] = 32'd61;
     memory[3592] = 32'd60;
     memory[3593] = 32'd242;
     memory[3594] = 32'd161;
     memory[3595] = 32'd54;
     memory[3596] = 32'd175;
     memory[3597] = 32'd192;
     memory[3598] = 32'd147;
     memory[3599] = 32'd210;
     memory[3600] = 32'd140;
     memory[3601] = 32'd198;
     memory[3602] = 32'd152;
     memory[3603] = 32'd196;
     memory[3604] = 32'd145;
     memory[3605] = 32'd59;
     memory[3606] = 32'd235;
     memory[3607] = 32'd36;
     memory[3608] = 32'd93;
     memory[3609] = 32'd59;
     memory[3610] = 32'd122;
     memory[3611] = 32'd68;
     memory[3612] = 32'd231;
     memory[3613] = 32'd250;
     memory[3614] = 32'd101;
     memory[3615] = 32'd100;
     memory[3616] = 32'd135;
     memory[3617] = 32'd56;
     memory[3618] = 32'd183;
     memory[3619] = 32'd246;
     memory[3620] = 32'd193;
     memory[3621] = 32'd206;
     memory[3622] = 32'd46;
     memory[3623] = 32'd127;
     memory[3624] = 32'd192;
     memory[3625] = 32'd200;
     memory[3626] = 32'd142;
     memory[3627] = 32'd118;
     memory[3628] = 32'd107;
     memory[3629] = 32'd149;
     memory[3630] = 32'd201;
     memory[3631] = 32'd93;
     memory[3632] = 32'd25;
     memory[3633] = 32'd71;
     memory[3634] = 32'd71;
     memory[3635] = 32'd93;
     memory[3636] = 32'd4;
     memory[3637] = 32'd157;
     memory[3638] = 32'd157;
     memory[3639] = 32'd242;
     memory[3640] = 32'd93;
     memory[3641] = 32'd77;
     memory[3642] = 32'd105;
     memory[3643] = 32'd86;
     memory[3644] = 32'd231;
     memory[3645] = 32'd81;
     memory[3646] = 32'd220;
     memory[3647] = 32'd75;
     memory[3648] = 32'd65;
     memory[3649] = 32'd161;
     memory[3650] = 32'd213;
     memory[3651] = 32'd166;
     memory[3652] = 32'd106;
     memory[3653] = 32'd130;
     memory[3654] = 32'd54;
     memory[3655] = 32'd230;
     memory[3656] = 32'd50;
     memory[3657] = 32'd101;
     memory[3658] = 32'd54;
     memory[3659] = 32'd228;
     memory[3660] = 32'd159;
     memory[3661] = 32'd31;
     memory[3662] = 32'd93;
     memory[3663] = 32'd55;
     memory[3664] = 32'd238;
     memory[3665] = 32'd242;
     memory[3666] = 32'd168;
     memory[3667] = 32'd91;
     memory[3668] = 32'd72;
     memory[3669] = 32'd205;
     memory[3670] = 32'd145;
     memory[3671] = 32'd246;
     memory[3672] = 32'd155;
     memory[3673] = 32'd32;
     memory[3674] = 32'd11;
     memory[3675] = 32'd107;
     memory[3676] = 32'd243;
     memory[3677] = 32'd92;
     memory[3678] = 32'd49;
     memory[3679] = 32'd208;
     memory[3680] = 32'd184;
     memory[3681] = 32'd110;
     memory[3682] = 32'd128;
     memory[3683] = 32'd112;
     memory[3684] = 32'd210;
     memory[3685] = 32'd215;
     memory[3686] = 32'd235;
     memory[3687] = 32'd198;
     memory[3688] = 32'd251;
     memory[3689] = 32'd54;
     memory[3690] = 32'd220;
     memory[3691] = 32'd173;
     memory[3692] = 32'd226;
     memory[3693] = 32'd124;
     memory[3694] = 32'd158;
     memory[3695] = 32'd115;
     memory[3696] = 32'd39;
     memory[3697] = 32'd92;
     memory[3698] = 32'd185;
     memory[3699] = 32'd99;
     memory[3700] = 32'd239;
     memory[3701] = 32'd182;
     memory[3702] = 32'd14;
     memory[3703] = 32'd230;
     memory[3704] = 32'd83;
     memory[3705] = 32'd206;
     memory[3706] = 32'd224;
     memory[3707] = 32'd54;
     memory[3708] = 32'd25;
     memory[3709] = 32'd53;
     memory[3710] = 32'd5;
     memory[3711] = 32'd100;
     memory[3712] = 32'd73;
     memory[3713] = 32'd181;
     memory[3714] = 32'd175;
     memory[3715] = 32'd44;
     memory[3716] = 32'd243;
     memory[3717] = 32'd196;
     memory[3718] = 32'd249;
     memory[3719] = 32'd176;
     memory[3720] = 32'd210;
     memory[3721] = 32'd167;
     memory[3722] = 32'd100;
     memory[3723] = 32'd13;
     memory[3724] = 32'd47;
     memory[3725] = 32'd223;
     memory[3726] = 32'd30;
     memory[3727] = 32'd142;
     memory[3728] = 32'd170;
     memory[3729] = 32'd200;
     memory[3730] = 32'd96;
     memory[3731] = 32'd157;
     memory[3732] = 32'd50;
     memory[3733] = 32'd162;
     memory[3734] = 32'd36;
     memory[3735] = 32'd56;
     memory[3736] = 32'd80;
     memory[3737] = 32'd109;
     memory[3738] = 32'd9;
     memory[3739] = 32'd190;
     memory[3740] = 32'd108;
     memory[3741] = 32'd140;
     memory[3742] = 32'd93;
     memory[3743] = 32'd172;
     memory[3744] = 32'd64;
     memory[3745] = 32'd152;
     memory[3746] = 32'd81;
     memory[3747] = 32'd134;
     memory[3748] = 32'd183;
     memory[3749] = 32'd138;
     memory[3750] = 32'd80;
     memory[3751] = 32'd12;
     memory[3752] = 32'd54;
     memory[3753] = 32'd197;
     memory[3754] = 32'd2;
     memory[3755] = 32'd2;
     memory[3756] = 32'd52;
     memory[3757] = 32'd209;
     memory[3758] = 32'd70;
     memory[3759] = 32'd0;
     memory[3760] = 32'd238;
     memory[3761] = 32'd249;
     memory[3762] = 32'd63;
     memory[3763] = 32'd75;
     memory[3764] = 32'd197;
     memory[3765] = 32'd251;
     memory[3766] = 32'd13;
     memory[3767] = 32'd137;
     memory[3768] = 32'd225;
     memory[3769] = 32'd99;
     memory[3770] = 32'd10;
     memory[3771] = 32'd212;
     memory[3772] = 32'd65;
     memory[3773] = 32'd2;
     memory[3774] = 32'd224;
     memory[3775] = 32'd150;
     memory[3776] = 32'd224;
     memory[3777] = 32'd15;
     memory[3778] = 32'd196;
     memory[3779] = 32'd106;
     memory[3780] = 32'd35;
     memory[3781] = 32'd187;
     memory[3782] = 32'd248;
     memory[3783] = 32'd246;
     memory[3784] = 32'd186;
     memory[3785] = 32'd193;
     memory[3786] = 32'd147;
     memory[3787] = 32'd74;
     memory[3788] = 32'd226;
     memory[3789] = 32'd160;
     memory[3790] = 32'd35;
     memory[3791] = 32'd77;
     memory[3792] = 32'd229;
     memory[3793] = 32'd239;
     memory[3794] = 32'd165;
     memory[3795] = 32'd82;
     memory[3796] = 32'd240;
     memory[3797] = 32'd108;
     memory[3798] = 32'd125;
     memory[3799] = 32'd192;
     memory[3800] = 32'd186;
     memory[3801] = 32'd177;
     memory[3802] = 32'd230;
     memory[3803] = 32'd137;
     memory[3804] = 32'd100;
     memory[3805] = 32'd88;
     memory[3806] = 32'd178;
     memory[3807] = 32'd182;
     memory[3808] = 32'd235;
     memory[3809] = 32'd148;
     memory[3810] = 32'd68;
     memory[3811] = 32'd67;
     memory[3812] = 32'd207;
     memory[3813] = 32'd9;
     memory[3814] = 32'd152;
     memory[3815] = 32'd175;
     memory[3816] = 32'd115;
     memory[3817] = 32'd216;
     memory[3818] = 32'd252;
     memory[3819] = 32'd188;
     memory[3820] = 32'd72;
     memory[3821] = 32'd2;
     memory[3822] = 32'd148;
     memory[3823] = 32'd32;
     memory[3824] = 32'd102;
     memory[3825] = 32'd115;
     memory[3826] = 32'd251;
     memory[3827] = 32'd157;
     memory[3828] = 32'd167;
     memory[3829] = 32'd219;
     memory[3830] = 32'd100;
     memory[3831] = 32'd208;
     memory[3832] = 32'd101;
     memory[3833] = 32'd78;
     memory[3834] = 32'd227;
     memory[3835] = 32'd52;
     memory[3836] = 32'd16;
     memory[3837] = 32'd247;
     memory[3838] = 32'd92;
     memory[3839] = 32'd83;
     memory[3840] = 32'd9;
     memory[3841] = 32'd22;
     memory[3842] = 32'd220;
     memory[3843] = 32'd56;
     memory[3844] = 32'd20;
     memory[3845] = 32'd13;
     memory[3846] = 32'd149;
     memory[3847] = 32'd158;
     memory[3848] = 32'd118;
     memory[3849] = 32'd197;
     memory[3850] = 32'd246;
     memory[3851] = 32'd185;
     memory[3852] = 32'd243;
     memory[3853] = 32'd209;
     memory[3854] = 32'd230;
     memory[3855] = 32'd72;
     memory[3856] = 32'd24;
     memory[3857] = 32'd26;
     memory[3858] = 32'd167;
     memory[3859] = 32'd66;
     memory[3860] = 32'd251;
     memory[3861] = 32'd216;
     memory[3862] = 32'd209;
     memory[3863] = 32'd30;
     memory[3864] = 32'd122;
     memory[3865] = 32'd123;
     memory[3866] = 32'd181;
     memory[3867] = 32'd29;
     memory[3868] = 32'd160;
     memory[3869] = 32'd93;
     memory[3870] = 32'd220;
     memory[3871] = 32'd179;
     memory[3872] = 32'd136;
     memory[3873] = 32'd93;
     memory[3874] = 32'd210;
     memory[3875] = 32'd200;
     memory[3876] = 32'd156;
     memory[3877] = 32'd190;
     memory[3878] = 32'd245;
     memory[3879] = 32'd95;
     memory[3880] = 32'd181;
     memory[3881] = 32'd215;
     memory[3882] = 32'd250;
     memory[3883] = 32'd138;
     memory[3884] = 32'd227;
     memory[3885] = 32'd19;
     memory[3886] = 32'd65;
     memory[3887] = 32'd133;
     memory[3888] = 32'd71;
     memory[3889] = 32'd237;
     memory[3890] = 32'd182;
     memory[3891] = 32'd236;
     memory[3892] = 32'd101;
     memory[3893] = 32'd114;
     memory[3894] = 32'd85;
     memory[3895] = 32'd241;
     memory[3896] = 32'd180;
     memory[3897] = 32'd151;
     memory[3898] = 32'd75;
     memory[3899] = 32'd93;
     memory[3900] = 32'd213;
     memory[3901] = 32'd244;
     memory[3902] = 32'd152;
     memory[3903] = 32'd52;
     memory[3904] = 32'd179;
     memory[3905] = 32'd201;
     memory[3906] = 32'd76;
     memory[3907] = 32'd124;
     memory[3908] = 32'd13;
     memory[3909] = 32'd204;
     memory[3910] = 32'd159;
     memory[3911] = 32'd249;
     memory[3912] = 32'd116;
     memory[3913] = 32'd171;
     memory[3914] = 32'd50;
     memory[3915] = 32'd117;
     memory[3916] = 32'd77;
     memory[3917] = 32'd122;
     memory[3918] = 32'd227;
     memory[3919] = 32'd50;
     memory[3920] = 32'd227;
     memory[3921] = 32'd96;
     memory[3922] = 32'd231;
     memory[3923] = 32'd120;
     memory[3924] = 32'd103;
     memory[3925] = 32'd56;
     memory[3926] = 32'd4;
     memory[3927] = 32'd57;
     memory[3928] = 32'd113;
     memory[3929] = 32'd232;
     memory[3930] = 32'd213;
     memory[3931] = 32'd94;
     memory[3932] = 32'd202;
     memory[3933] = 32'd210;
     memory[3934] = 32'd14;
     memory[3935] = 32'd142;
     memory[3936] = 32'd247;
     memory[3937] = 32'd56;
     memory[3938] = 32'd6;
     memory[3939] = 32'd204;
     memory[3940] = 32'd109;
     memory[3941] = 32'd212;
     memory[3942] = 32'd79;
     memory[3943] = 32'd18;
     memory[3944] = 32'd142;
     memory[3945] = 32'd223;
     memory[3946] = 32'd4;
     memory[3947] = 32'd223;
     memory[3948] = 32'd7;
     memory[3949] = 32'd250;
     memory[3950] = 32'd215;
     memory[3951] = 32'd123;
     memory[3952] = 32'd164;
     memory[3953] = 32'd75;
     memory[3954] = 32'd226;
     memory[3955] = 32'd117;
     memory[3956] = 32'd208;
     memory[3957] = 32'd126;
     memory[3958] = 32'd64;
     memory[3959] = 32'd131;
     memory[3960] = 32'd150;
     memory[3961] = 32'd239;
     memory[3962] = 32'd153;
     memory[3963] = 32'd145;
     memory[3964] = 32'd137;
     memory[3965] = 32'd56;
     memory[3966] = 32'd226;
     memory[3967] = 32'd155;
     memory[3968] = 32'd227;
     memory[3969] = 32'd166;
     memory[3970] = 32'd221;
     memory[3971] = 32'd22;
     memory[3972] = 32'd120;
     memory[3973] = 32'd44;
     memory[3974] = 32'd126;
     memory[3975] = 32'd252;
     memory[3976] = 32'd155;
     memory[3977] = 32'd251;
     memory[3978] = 32'd188;
     memory[3979] = 32'd203;
     memory[3980] = 32'd99;
     memory[3981] = 32'd82;
     memory[3982] = 32'd52;
     memory[3983] = 32'd68;
     memory[3984] = 32'd171;
     memory[3985] = 32'd63;
     memory[3986] = 32'd202;
     memory[3987] = 32'd109;
     memory[3988] = 32'd83;
     memory[3989] = 32'd79;
     memory[3990] = 32'd180;
     memory[3991] = 32'd144;
     memory[3992] = 32'd67;
     memory[3993] = 32'd38;
     memory[3994] = 32'd97;
     memory[3995] = 32'd73;
     memory[3996] = 32'd168;
     memory[3997] = 32'd249;
     memory[3998] = 32'd83;
     memory[3999] = 32'd20;
     memory[4000] = 32'd0;
     memory[4001] = 32'd95;
     memory[4002] = 32'd254;
     memory[4003] = 32'd19;
     memory[4004] = 32'd196;
     memory[4005] = 32'd88;
     memory[4006] = 32'd96;
     memory[4007] = 32'd29;
     memory[4008] = 32'd77;
     memory[4009] = 32'd236;
     memory[4010] = 32'd32;
     memory[4011] = 32'd127;
     memory[4012] = 32'd118;
     memory[4013] = 32'd140;
     memory[4014] = 32'd68;
     memory[4015] = 32'd111;
     memory[4016] = 32'd175;
     memory[4017] = 32'd232;
     memory[4018] = 32'd81;
     memory[4019] = 32'd137;
     memory[4020] = 32'd240;
     memory[4021] = 32'd150;
     memory[4022] = 32'd97;
     memory[4023] = 32'd221;
     memory[4024] = 32'd35;
     memory[4025] = 32'd239;
     memory[4026] = 32'd216;
     memory[4027] = 32'd87;
     memory[4028] = 32'd149;
     memory[4029] = 32'd87;
     memory[4030] = 32'd189;
     memory[4031] = 32'd215;
     memory[4032] = 32'd239;
     memory[4033] = 32'd25;
     memory[4034] = 32'd122;
     memory[4035] = 32'd3;
     memory[4036] = 32'd94;
     memory[4037] = 32'd132;
     memory[4038] = 32'd196;
     memory[4039] = 32'd9;
     memory[4040] = 32'd235;
     memory[4041] = 32'd75;
     memory[4042] = 32'd83;
     memory[4043] = 32'd240;
     memory[4044] = 32'd137;
     memory[4045] = 32'd204;
     memory[4046] = 32'd248;
     memory[4047] = 32'd149;
     memory[4048] = 32'd193;
     memory[4049] = 32'd185;
     memory[4050] = 32'd194;
     memory[4051] = 32'd183;
     memory[4052] = 32'd53;
     memory[4053] = 32'd225;
     memory[4054] = 32'd157;
     memory[4055] = 32'd204;
     memory[4056] = 32'd223;
     memory[4057] = 32'd95;
     memory[4058] = 32'd15;
     memory[4059] = 32'd239;
     memory[4060] = 32'd228;
     memory[4061] = 32'd81;
     memory[4062] = 32'd31;
     memory[4063] = 32'd122;
     memory[4064] = 32'd67;
     memory[4065] = 32'd133;
     memory[4066] = 32'd89;
     memory[4067] = 32'd188;
     memory[4068] = 32'd146;
     memory[4069] = 32'd30;
     memory[4070] = 32'd191;
     memory[4071] = 32'd248;
     memory[4072] = 32'd9;
     memory[4073] = 32'd179;
     memory[4074] = 32'd21;
     memory[4075] = 32'd97;
     memory[4076] = 32'd243;
     memory[4077] = 32'd239;
     memory[4078] = 32'd139;
     memory[4079] = 32'd180;
     memory[4080] = 32'd243;
     memory[4081] = 32'd117;
     memory[4082] = 32'd24;
     memory[4083] = 32'd119;
     memory[4084] = 32'd110;
     memory[4085] = 32'd8;
     memory[4086] = 32'd241;
     memory[4087] = 32'd45;
     memory[4088] = 32'd41;
     memory[4089] = 32'd58;
     memory[4090] = 32'd177;
     memory[4091] = 32'd219;
     memory[4092] = 32'd223;
     memory[4093] = 32'd207;
     memory[4094] = 32'd158;
     memory[4095] = 32'd159;
     memory[4096] = 32'd247;
     memory[4097] = 32'd28;   //begining of matrix B
     memory[4098] = 32'd81;
     memory[4099] = 32'd57;
     memory[4100] = 32'd16;
     memory[4101] = 32'd27;
     memory[4102] = 32'd28;
     memory[4103] = 32'd38;
     memory[4104] = 32'd26;
     memory[4105] = 32'd17;
     memory[4106] = 32'd51;
     memory[4107] = 32'd62;
     memory[4108] = 32'd18;
     memory[4109] = 32'd35;
     memory[4110] = 32'd19;
     memory[4111] = 32'd10;
     memory[4112] = 32'd73;
     memory[4113] = 32'd100;
     memory[4114] = 32'd208;
     memory[4115] = 32'd124;
     memory[4116] = 32'd194;
     memory[4117] = 32'd187;
     memory[4118] = 32'd11;
     memory[4119] = 32'd221;
     memory[4120] = 32'd205;
     memory[4121] = 32'd129;
     memory[4122] = 32'd164;
     memory[4123] = 32'd182;
     memory[4124] = 32'd142;
     memory[4125] = 32'd113;
     memory[4126] = 32'd72;
     memory[4127] = 32'd199;
     memory[4128] = 32'd86;
     memory[4129] = 32'd31;
     memory[4130] = 32'd150;
     memory[4131] = 32'd251;
     memory[4132] = 32'd150;
     memory[4133] = 32'd85;
     memory[4134] = 32'd25;
     memory[4135] = 32'd20;
     memory[4136] = 32'd89;
     memory[4137] = 32'd248;
     memory[4138] = 32'd189;
     memory[4139] = 32'd35;
     memory[4140] = 32'd181;
     memory[4141] = 32'd201;
     memory[4142] = 32'd212;
     memory[4143] = 32'd207;
     memory[4144] = 32'd13;
     memory[4145] = 32'd95;
     memory[4146] = 32'd167;
     memory[4147] = 32'd46;
     memory[4148] = 32'd84;
     memory[4149] = 32'd225;
     memory[4150] = 32'd89;
     memory[4151] = 32'd181;
     memory[4152] = 32'd168;
     memory[4153] = 32'd98;
     memory[4154] = 32'd72;
     memory[4155] = 32'd58;
     memory[4156] = 32'd42;
     memory[4157] = 32'd163;
     memory[4158] = 32'd83;
     memory[4159] = 32'd15;
     memory[4160] = 32'd157;
     memory[4161] = 32'd248;
     memory[4162] = 32'd179;
     memory[4163] = 32'd210;
     memory[4164] = 32'd208;
     memory[4165] = 32'd122;
     memory[4166] = 32'd206;
     memory[4167] = 32'd11;
     memory[4168] = 32'd121;
     memory[4169] = 32'd189;
     memory[4170] = 32'd56;
     memory[4171] = 32'd123;
     memory[4172] = 32'd19;
     memory[4173] = 32'd113;
     memory[4174] = 32'd160;
     memory[4175] = 32'd185;
     memory[4176] = 32'd190;
     memory[4177] = 32'd8;
     memory[4178] = 32'd39;
     memory[4179] = 32'd111;
     memory[4180] = 32'd212;
     memory[4181] = 32'd57;
     memory[4182] = 32'd161;
     memory[4183] = 32'd219;
     memory[4184] = 32'd3;
     memory[4185] = 32'd233;
     memory[4186] = 32'd15;
     memory[4187] = 32'd38;
     memory[4188] = 32'd198;
     memory[4189] = 32'd80;
     memory[4190] = 32'd232;
     memory[4191] = 32'd193;
     memory[4192] = 32'd89;
     memory[4193] = 32'd39;
     memory[4194] = 32'd167;
     memory[4195] = 32'd20;
     memory[4196] = 32'd238;
     memory[4197] = 32'd41;
     memory[4198] = 32'd54;
     memory[4199] = 32'd71;
     memory[4200] = 32'd92;
     memory[4201] = 32'd122;
     memory[4202] = 32'd45;
     memory[4203] = 32'd210;
     memory[4204] = 32'd254;
     memory[4205] = 32'd74;
     memory[4206] = 32'd40;
     memory[4207] = 32'd85;
     memory[4208] = 32'd226;
     memory[4209] = 32'd170;
     memory[4210] = 32'd113;
     memory[4211] = 32'd253;
     memory[4212] = 32'd230;
     memory[4213] = 32'd196;
     memory[4214] = 32'd122;
     memory[4215] = 32'd68;
     memory[4216] = 32'd128;
     memory[4217] = 32'd84;
     memory[4218] = 32'd219;
     memory[4219] = 32'd217;
     memory[4220] = 32'd27;
     memory[4221] = 32'd50;
     memory[4222] = 32'd123;
     memory[4223] = 32'd70;
     memory[4224] = 32'd198;
     memory[4225] = 32'd250;
     memory[4226] = 32'd195;
     memory[4227] = 32'd40;
     memory[4228] = 32'd189;
     memory[4229] = 32'd137;
     memory[4230] = 32'd31;
     memory[4231] = 32'd75;
     memory[4232] = 32'd163;
     memory[4233] = 32'd134;
     memory[4234] = 32'd173;
     memory[4235] = 32'd89;
     memory[4236] = 32'd139;
     memory[4237] = 32'd190;
     memory[4238] = 32'd103;
     memory[4239] = 32'd177;
     memory[4240] = 32'd121;
     memory[4241] = 32'd114;
     memory[4242] = 32'd239;
     memory[4243] = 32'd46;
     memory[4244] = 32'd67;
     memory[4245] = 32'd199;
     memory[4246] = 32'd115;
     memory[4247] = 32'd81;
     memory[4248] = 32'd54;
     memory[4249] = 32'd52;
     memory[4250] = 32'd148;
     memory[4251] = 32'd32;
     memory[4252] = 32'd109;
     memory[4253] = 32'd151;
     memory[4254] = 32'd179;
     memory[4255] = 32'd20;
     memory[4256] = 32'd135;
     memory[4257] = 32'd172;
     memory[4258] = 32'd66;
     memory[4259] = 32'd84;
     memory[4260] = 32'd224;
     memory[4261] = 32'd96;
     memory[4262] = 32'd13;
     memory[4263] = 32'd242;
     memory[4264] = 32'd251;
     memory[4265] = 32'd3;
     memory[4266] = 32'd138;
     memory[4267] = 32'd240;
     memory[4268] = 32'd0;
     memory[4269] = 32'd170;
     memory[4270] = 32'd105;
     memory[4271] = 32'd229;
     memory[4272] = 32'd94;
     memory[4273] = 32'd245;
     memory[4274] = 32'd222;
     memory[4275] = 32'd150;
     memory[4276] = 32'd21;
     memory[4277] = 32'd33;
     memory[4278] = 32'd110;
     memory[4279] = 32'd21;
     memory[4280] = 32'd82;
     memory[4281] = 32'd191;
     memory[4282] = 32'd47;
     memory[4283] = 32'd159;
     memory[4284] = 32'd85;
     memory[4285] = 32'd6;
     memory[4286] = 32'd140;
     memory[4287] = 32'd90;
     memory[4288] = 32'd136;
     memory[4289] = 32'd155;
     memory[4290] = 32'd106;
     memory[4291] = 32'd222;
     memory[4292] = 32'd18;
     memory[4293] = 32'd122;
     memory[4294] = 32'd64;
     memory[4295] = 32'd26;
     memory[4296] = 32'd62;
     memory[4297] = 32'd231;
     memory[4298] = 32'd157;
     memory[4299] = 32'd8;
     memory[4300] = 32'd201;
     memory[4301] = 32'd77;
     memory[4302] = 32'd221;
     memory[4303] = 32'd17;
     memory[4304] = 32'd75;
     memory[4305] = 32'd44;
     memory[4306] = 32'd201;
     memory[4307] = 32'd137;
     memory[4308] = 32'd4;
     memory[4309] = 32'd91;
     memory[4310] = 32'd220;
     memory[4311] = 32'd172;
     memory[4312] = 32'd32;
     memory[4313] = 32'd96;
     memory[4314] = 32'd33;
     memory[4315] = 32'd71;
     memory[4316] = 32'd219;
     memory[4317] = 32'd78;
     memory[4318] = 32'd94;
     memory[4319] = 32'd125;
     memory[4320] = 32'd132;
     memory[4321] = 32'd32;
     memory[4322] = 32'd78;
     memory[4323] = 32'd124;
     memory[4324] = 32'd75;
     memory[4325] = 32'd107;
     memory[4326] = 32'd80;
     memory[4327] = 32'd58;
     memory[4328] = 32'd117;
     memory[4329] = 32'd64;
     memory[4330] = 32'd166;
     memory[4331] = 32'd204;
     memory[4332] = 32'd74;
     memory[4333] = 32'd79;
     memory[4334] = 32'd216;
     memory[4335] = 32'd218;
     memory[4336] = 32'd218;
     memory[4337] = 32'd75;
     memory[4338] = 32'd30;
     memory[4339] = 32'd201;
     memory[4340] = 32'd98;
     memory[4341] = 32'd94;
     memory[4342] = 32'd38;
     memory[4343] = 32'd208;
     memory[4344] = 32'd233;
     memory[4345] = 32'd238;
     memory[4346] = 32'd154;
     memory[4347] = 32'd188;
     memory[4348] = 32'd76;
     memory[4349] = 32'd178;
     memory[4350] = 32'd124;
     memory[4351] = 32'd8;
     memory[4352] = 32'd59;
     memory[4353] = 32'd160;
     memory[4354] = 32'd184;
     memory[4355] = 32'd50;
     memory[4356] = 32'd251;
     memory[4357] = 32'd187;
     memory[4358] = 32'd59;
     memory[4359] = 32'd139;
     memory[4360] = 32'd109;
     memory[4361] = 32'd252;
     memory[4362] = 32'd73;
     memory[4363] = 32'd145;
     memory[4364] = 32'd113;
     memory[4365] = 32'd182;
     memory[4366] = 32'd237;
     memory[4367] = 32'd149;
     memory[4368] = 32'd187;
     memory[4369] = 32'd105;
     memory[4370] = 32'd211;
     memory[4371] = 32'd86;
     memory[4372] = 32'd60;
     memory[4373] = 32'd122;
     memory[4374] = 32'd114;
     memory[4375] = 32'd16;
     memory[4376] = 32'd174;
     memory[4377] = 32'd126;
     memory[4378] = 32'd144;
     memory[4379] = 32'd3;
     memory[4380] = 32'd114;
     memory[4381] = 32'd101;
     memory[4382] = 32'd135;
     memory[4383] = 32'd17;
     memory[4384] = 32'd252;
     memory[4385] = 32'd93;
     memory[4386] = 32'd57;
     memory[4387] = 32'd250;
     memory[4388] = 32'd26;
     memory[4389] = 32'd56;
     memory[4390] = 32'd168;
     memory[4391] = 32'd197;
     memory[4392] = 32'd34;
     memory[4393] = 32'd179;
     memory[4394] = 32'd71;
     memory[4395] = 32'd26;
     memory[4396] = 32'd123;
     memory[4397] = 32'd94;
     memory[4398] = 32'd14;
     memory[4399] = 32'd238;
     memory[4400] = 32'd86;
     memory[4401] = 32'd33;
     memory[4402] = 32'd184;
     memory[4403] = 32'd58;
     memory[4404] = 32'd121;
     memory[4405] = 32'd183;
     memory[4406] = 32'd49;
     memory[4407] = 32'd107;
     memory[4408] = 32'd63;
     memory[4409] = 32'd125;
     memory[4410] = 32'd145;
     memory[4411] = 32'd102;
     memory[4412] = 32'd224;
     memory[4413] = 32'd246;
     memory[4414] = 32'd91;
     memory[4415] = 32'd172;
     memory[4416] = 32'd156;
     memory[4417] = 32'd229;
     memory[4418] = 32'd130;
     memory[4419] = 32'd167;
     memory[4420] = 32'd25;
     memory[4421] = 32'd139;
     memory[4422] = 32'd195;
     memory[4423] = 32'd97;
     memory[4424] = 32'd116;
     memory[4425] = 32'd62;
     memory[4426] = 32'd25;
     memory[4427] = 32'd220;
     memory[4428] = 32'd65;
     memory[4429] = 32'd239;
     memory[4430] = 32'd184;
     memory[4431] = 32'd89;
     memory[4432] = 32'd26;
     memory[4433] = 32'd5;
     memory[4434] = 32'd152;
     memory[4435] = 32'd250;
     memory[4436] = 32'd245;
     memory[4437] = 32'd121;
     memory[4438] = 32'd180;
     memory[4439] = 32'd83;
     memory[4440] = 32'd108;
     memory[4441] = 32'd107;
     memory[4442] = 32'd135;
     memory[4443] = 32'd207;
     memory[4444] = 32'd26;
     memory[4445] = 32'd194;
     memory[4446] = 32'd12;
     memory[4447] = 32'd219;
     memory[4448] = 32'd251;
     memory[4449] = 32'd153;
     memory[4450] = 32'd106;
     memory[4451] = 32'd28;
     memory[4452] = 32'd83;
     memory[4453] = 32'd110;
     memory[4454] = 32'd254;
     memory[4455] = 32'd251;
     memory[4456] = 32'd57;
     memory[4457] = 32'd54;
     memory[4458] = 32'd80;
     memory[4459] = 32'd18;
     memory[4460] = 32'd236;
     memory[4461] = 32'd122;
     memory[4462] = 32'd179;
     memory[4463] = 32'd245;
     memory[4464] = 32'd249;
     memory[4465] = 32'd47;
     memory[4466] = 32'd3;
     memory[4467] = 32'd49;
     memory[4468] = 32'd22;
     memory[4469] = 32'd199;
     memory[4470] = 32'd42;
     memory[4471] = 32'd55;
     memory[4472] = 32'd21;
     memory[4473] = 32'd102;
     memory[4474] = 32'd209;
     memory[4475] = 32'd118;
     memory[4476] = 32'd103;
     memory[4477] = 32'd214;
     memory[4478] = 32'd245;
     memory[4479] = 32'd155;
     memory[4480] = 32'd110;
     memory[4481] = 32'd31;
     memory[4482] = 32'd91;
     memory[4483] = 32'd27;
     memory[4484] = 32'd105;
     memory[4485] = 32'd206;
     memory[4486] = 32'd235;
     memory[4487] = 32'd52;
     memory[4488] = 32'd199;
     memory[4489] = 32'd116;
     memory[4490] = 32'd115;
     memory[4491] = 32'd44;
     memory[4492] = 32'd200;
     memory[4493] = 32'd0;
     memory[4494] = 32'd176;
     memory[4495] = 32'd59;
     memory[4496] = 32'd10;
     memory[4497] = 32'd34;
     memory[4498] = 32'd48;
     memory[4499] = 32'd192;
     memory[4500] = 32'd61;
     memory[4501] = 32'd220;
     memory[4502] = 32'd189;
     memory[4503] = 32'd242;
     memory[4504] = 32'd56;
     memory[4505] = 32'd23;
     memory[4506] = 32'd151;
     memory[4507] = 32'd197;
     memory[4508] = 32'd105;
     memory[4509] = 32'd35;
     memory[4510] = 32'd127;
     memory[4511] = 32'd87;
     memory[4512] = 32'd197;
     memory[4513] = 32'd188;
     memory[4514] = 32'd1;
     memory[4515] = 32'd74;
     memory[4516] = 32'd159;
     memory[4517] = 32'd228;
     memory[4518] = 32'd35;
     memory[4519] = 32'd57;
     memory[4520] = 32'd135;
     memory[4521] = 32'd197;
     memory[4522] = 32'd11;
     memory[4523] = 32'd3;
     memory[4524] = 32'd157;
     memory[4525] = 32'd28;
     memory[4526] = 32'd123;
     memory[4527] = 32'd101;
     memory[4528] = 32'd1;
     memory[4529] = 32'd4;
     memory[4530] = 32'd43;
     memory[4531] = 32'd200;
     memory[4532] = 32'd248;
     memory[4533] = 32'd150;
     memory[4534] = 32'd24;
     memory[4535] = 32'd185;
     memory[4536] = 32'd247;
     memory[4537] = 32'd25;
     memory[4538] = 32'd69;
     memory[4539] = 32'd33;
     memory[4540] = 32'd49;
     memory[4541] = 32'd94;
     memory[4542] = 32'd186;
     memory[4543] = 32'd236;
     memory[4544] = 32'd144;
     memory[4545] = 32'd84;
     memory[4546] = 32'd199;
     memory[4547] = 32'd106;
     memory[4548] = 32'd225;
     memory[4549] = 32'd198;
     memory[4550] = 32'd98;
     memory[4551] = 32'd65;
     memory[4552] = 32'd247;
     memory[4553] = 32'd179;
     memory[4554] = 32'd79;
     memory[4555] = 32'd132;
     memory[4556] = 32'd222;
     memory[4557] = 32'd99;
     memory[4558] = 32'd38;
     memory[4559] = 32'd158;
     memory[4560] = 32'd210;
     memory[4561] = 32'd158;
     memory[4562] = 32'd170;
     memory[4563] = 32'd144;
     memory[4564] = 32'd226;
     memory[4565] = 32'd175;
     memory[4566] = 32'd15;
     memory[4567] = 32'd131;
     memory[4568] = 32'd2;
     memory[4569] = 32'd170;
     memory[4570] = 32'd83;
     memory[4571] = 32'd238;
     memory[4572] = 32'd5;
     memory[4573] = 32'd129;
     memory[4574] = 32'd176;
     memory[4575] = 32'd171;
     memory[4576] = 32'd202;
     memory[4577] = 32'd35;
     memory[4578] = 32'd244;
     memory[4579] = 32'd220;
     memory[4580] = 32'd207;
     memory[4581] = 32'd62;
     memory[4582] = 32'd231;
     memory[4583] = 32'd98;
     memory[4584] = 32'd240;
     memory[4585] = 32'd199;
     memory[4586] = 32'd234;
     memory[4587] = 32'd208;
     memory[4588] = 32'd125;
     memory[4589] = 32'd162;
     memory[4590] = 32'd148;
     memory[4591] = 32'd225;
     memory[4592] = 32'd36;
     memory[4593] = 32'd239;
     memory[4594] = 32'd59;
     memory[4595] = 32'd172;
     memory[4596] = 32'd34;
     memory[4597] = 32'd37;
     memory[4598] = 32'd19;
     memory[4599] = 32'd78;
     memory[4600] = 32'd190;
     memory[4601] = 32'd230;
     memory[4602] = 32'd132;
     memory[4603] = 32'd190;
     memory[4604] = 32'd132;
     memory[4605] = 32'd117;
     memory[4606] = 32'd15;
     memory[4607] = 32'd14;
     memory[4608] = 32'd39;
     memory[4609] = 32'd155;
     memory[4610] = 32'd181;
     memory[4611] = 32'd120;
     memory[4612] = 32'd111;
     memory[4613] = 32'd231;
     memory[4614] = 32'd52;
     memory[4615] = 32'd180;
     memory[4616] = 32'd77;
     memory[4617] = 32'd16;
     memory[4618] = 32'd55;
     memory[4619] = 32'd38;
     memory[4620] = 32'd150;
     memory[4621] = 32'd51;
     memory[4622] = 32'd188;
     memory[4623] = 32'd48;
     memory[4624] = 32'd77;
     memory[4625] = 32'd8;
     memory[4626] = 32'd248;
     memory[4627] = 32'd139;
     memory[4628] = 32'd92;
     memory[4629] = 32'd173;
     memory[4630] = 32'd5;
     memory[4631] = 32'd114;
     memory[4632] = 32'd46;
     memory[4633] = 32'd145;
     memory[4634] = 32'd139;
     memory[4635] = 32'd52;
     memory[4636] = 32'd195;
     memory[4637] = 32'd50;
     memory[4638] = 32'd248;
     memory[4639] = 32'd25;
     memory[4640] = 32'd10;
     memory[4641] = 32'd61;
     memory[4642] = 32'd136;
     memory[4643] = 32'd196;
     memory[4644] = 32'd78;
     memory[4645] = 32'd148;
     memory[4646] = 32'd98;
     memory[4647] = 32'd216;
     memory[4648] = 32'd83;
     memory[4649] = 32'd242;
     memory[4650] = 32'd216;
     memory[4651] = 32'd111;
     memory[4652] = 32'd253;
     memory[4653] = 32'd14;
     memory[4654] = 32'd22;
     memory[4655] = 32'd47;
     memory[4656] = 32'd14;
     memory[4657] = 32'd201;
     memory[4658] = 32'd251;
     memory[4659] = 32'd27;
     memory[4660] = 32'd45;
     memory[4661] = 32'd10;
     memory[4662] = 32'd215;
     memory[4663] = 32'd206;
     memory[4664] = 32'd194;
     memory[4665] = 32'd23;
     memory[4666] = 32'd2;
     memory[4667] = 32'd253;
     memory[4668] = 32'd130;
     memory[4669] = 32'd59;
     memory[4670] = 32'd66;
     memory[4671] = 32'd213;
     memory[4672] = 32'd251;
     memory[4673] = 32'd91;
     memory[4674] = 32'd105;
     memory[4675] = 32'd70;
     memory[4676] = 32'd112;
     memory[4677] = 32'd254;
     memory[4678] = 32'd236;
     memory[4679] = 32'd161;
     memory[4680] = 32'd155;
     memory[4681] = 32'd102;
     memory[4682] = 32'd224;
     memory[4683] = 32'd9;
     memory[4684] = 32'd114;
     memory[4685] = 32'd205;
     memory[4686] = 32'd88;
     memory[4687] = 32'd88;
     memory[4688] = 32'd63;
     memory[4689] = 32'd219;
     memory[4690] = 32'd84;
     memory[4691] = 32'd168;
     memory[4692] = 32'd118;
     memory[4693] = 32'd149;
     memory[4694] = 32'd211;
     memory[4695] = 32'd18;
     memory[4696] = 32'd250;
     memory[4697] = 32'd157;
     memory[4698] = 32'd52;
     memory[4699] = 32'd89;
     memory[4700] = 32'd28;
     memory[4701] = 32'd91;
     memory[4702] = 32'd8;
     memory[4703] = 32'd209;
     memory[4704] = 32'd75;
     memory[4705] = 32'd173;
     memory[4706] = 32'd51;
     memory[4707] = 32'd153;
     memory[4708] = 32'd161;
     memory[4709] = 32'd0;
     memory[4710] = 32'd20;
     memory[4711] = 32'd184;
     memory[4712] = 32'd54;
     memory[4713] = 32'd179;
     memory[4714] = 32'd207;
     memory[4715] = 32'd22;
     memory[4716] = 32'd185;
     memory[4717] = 32'd137;
     memory[4718] = 32'd67;
     memory[4719] = 32'd63;
     memory[4720] = 32'd14;
     memory[4721] = 32'd172;
     memory[4722] = 32'd165;
     memory[4723] = 32'd102;
     memory[4724] = 32'd224;
     memory[4725] = 32'd225;
     memory[4726] = 32'd48;
     memory[4727] = 32'd220;
     memory[4728] = 32'd208;
     memory[4729] = 32'd29;
     memory[4730] = 32'd120;
     memory[4731] = 32'd3;
     memory[4732] = 32'd34;
     memory[4733] = 32'd116;
     memory[4734] = 32'd224;
     memory[4735] = 32'd22;
     memory[4736] = 32'd242;
     memory[4737] = 32'd49;
     memory[4738] = 32'd251;
     memory[4739] = 32'd184;
     memory[4740] = 32'd30;
     memory[4741] = 32'd166;
     memory[4742] = 32'd68;
     memory[4743] = 32'd30;
     memory[4744] = 32'd59;
     memory[4745] = 32'd32;
     memory[4746] = 32'd3;
     memory[4747] = 32'd48;
     memory[4748] = 32'd3;
     memory[4749] = 32'd173;
     memory[4750] = 32'd198;
     memory[4751] = 32'd32;
     memory[4752] = 32'd111;
     memory[4753] = 32'd183;
     memory[4754] = 32'd108;
     memory[4755] = 32'd116;
     memory[4756] = 32'd168;
     memory[4757] = 32'd177;
     memory[4758] = 32'd14;
     memory[4759] = 32'd0;
     memory[4760] = 32'd148;
     memory[4761] = 32'd72;
     memory[4762] = 32'd68;
     memory[4763] = 32'd105;
     memory[4764] = 32'd92;
     memory[4765] = 32'd235;
     memory[4766] = 32'd81;
     memory[4767] = 32'd76;
     memory[4768] = 32'd57;
     memory[4769] = 32'd114;
     memory[4770] = 32'd244;
     memory[4771] = 32'd159;
     memory[4772] = 32'd23;
     memory[4773] = 32'd79;
     memory[4774] = 32'd104;
     memory[4775] = 32'd79;
     memory[4776] = 32'd129;
     memory[4777] = 32'd83;
     memory[4778] = 32'd188;
     memory[4779] = 32'd61;
     memory[4780] = 32'd18;
     memory[4781] = 32'd247;
     memory[4782] = 32'd135;
     memory[4783] = 32'd245;
     memory[4784] = 32'd141;
     memory[4785] = 32'd180;
     memory[4786] = 32'd105;
     memory[4787] = 32'd130;
     memory[4788] = 32'd21;
     memory[4789] = 32'd86;
     memory[4790] = 32'd25;
     memory[4791] = 32'd78;
     memory[4792] = 32'd147;
     memory[4793] = 32'd201;
     memory[4794] = 32'd91;
     memory[4795] = 32'd249;
     memory[4796] = 32'd182;
     memory[4797] = 32'd249;
     memory[4798] = 32'd249;
     memory[4799] = 32'd77;
     memory[4800] = 32'd88;
     memory[4801] = 32'd200;
     memory[4802] = 32'd161;
     memory[4803] = 32'd252;
     memory[4804] = 32'd115;
     memory[4805] = 32'd239;
     memory[4806] = 32'd1;
     memory[4807] = 32'd59;
     memory[4808] = 32'd176;
     memory[4809] = 32'd77;
     memory[4810] = 32'd193;
     memory[4811] = 32'd96;
     memory[4812] = 32'd152;
     memory[4813] = 32'd79;
     memory[4814] = 32'd88;
     memory[4815] = 32'd174;
     memory[4816] = 32'd169;
     memory[4817] = 32'd66;
     memory[4818] = 32'd140;
     memory[4819] = 32'd56;
     memory[4820] = 32'd10;
     memory[4821] = 32'd223;
     memory[4822] = 32'd250;
     memory[4823] = 32'd38;
     memory[4824] = 32'd189;
     memory[4825] = 32'd21;
     memory[4826] = 32'd19;
     memory[4827] = 32'd217;
     memory[4828] = 32'd2;
     memory[4829] = 32'd119;
     memory[4830] = 32'd174;
     memory[4831] = 32'd68;
     memory[4832] = 32'd40;
     memory[4833] = 32'd84;
     memory[4834] = 32'd102;
     memory[4835] = 32'd175;
     memory[4836] = 32'd120;
     memory[4837] = 32'd63;
     memory[4838] = 32'd78;
     memory[4839] = 32'd188;
     memory[4840] = 32'd226;
     memory[4841] = 32'd214;
     memory[4842] = 32'd98;
     memory[4843] = 32'd1;
     memory[4844] = 32'd82;
     memory[4845] = 32'd218;
     memory[4846] = 32'd63;
     memory[4847] = 32'd39;
     memory[4848] = 32'd170;
     memory[4849] = 32'd138;
     memory[4850] = 32'd187;
     memory[4851] = 32'd19;
     memory[4852] = 32'd128;
     memory[4853] = 32'd134;
     memory[4854] = 32'd126;
     memory[4855] = 32'd185;
     memory[4856] = 32'd116;
     memory[4857] = 32'd141;
     memory[4858] = 32'd30;
     memory[4859] = 32'd208;
     memory[4860] = 32'd55;
     memory[4861] = 32'd241;
     memory[4862] = 32'd233;
     memory[4863] = 32'd50;
     memory[4864] = 32'd242;
     memory[4865] = 32'd134;
     memory[4866] = 32'd253;
     memory[4867] = 32'd210;
     memory[4868] = 32'd207;
     memory[4869] = 32'd208;
     memory[4870] = 32'd136;
     memory[4871] = 32'd9;
     memory[4872] = 32'd28;
     memory[4873] = 32'd132;
     memory[4874] = 32'd89;
     memory[4875] = 32'd34;
     memory[4876] = 32'd56;
     memory[4877] = 32'd180;
     memory[4878] = 32'd67;
     memory[4879] = 32'd124;
     memory[4880] = 32'd69;
     memory[4881] = 32'd22;
     memory[4882] = 32'd188;
     memory[4883] = 32'd143;
     memory[4884] = 32'd56;
     memory[4885] = 32'd144;
     memory[4886] = 32'd175;
     memory[4887] = 32'd192;
     memory[4888] = 32'd64;
     memory[4889] = 32'd119;
     memory[4890] = 32'd129;
     memory[4891] = 32'd5;
     memory[4892] = 32'd179;
     memory[4893] = 32'd58;
     memory[4894] = 32'd83;
     memory[4895] = 32'd67;
     memory[4896] = 32'd30;
     memory[4897] = 32'd61;
     memory[4898] = 32'd68;
     memory[4899] = 32'd33;
     memory[4900] = 32'd249;
     memory[4901] = 32'd157;
     memory[4902] = 32'd143;
     memory[4903] = 32'd200;
     memory[4904] = 32'd209;
     memory[4905] = 32'd228;
     memory[4906] = 32'd197;
     memory[4907] = 32'd17;
     memory[4908] = 32'd146;
     memory[4909] = 32'd65;
     memory[4910] = 32'd254;
     memory[4911] = 32'd86;
     memory[4912] = 32'd6;
     memory[4913] = 32'd174;
     memory[4914] = 32'd157;
     memory[4915] = 32'd18;
     memory[4916] = 32'd203;
     memory[4917] = 32'd248;
     memory[4918] = 32'd32;
     memory[4919] = 32'd208;
     memory[4920] = 32'd182;
     memory[4921] = 32'd154;
     memory[4922] = 32'd87;
     memory[4923] = 32'd173;
     memory[4924] = 32'd144;
     memory[4925] = 32'd223;
     memory[4926] = 32'd4;
     memory[4927] = 32'd186;
     memory[4928] = 32'd180;
     memory[4929] = 32'd166;
     memory[4930] = 32'd201;
     memory[4931] = 32'd114;
     memory[4932] = 32'd100;
     memory[4933] = 32'd30;
     memory[4934] = 32'd136;
     memory[4935] = 32'd143;
     memory[4936] = 32'd233;
     memory[4937] = 32'd86;
     memory[4938] = 32'd82;
     memory[4939] = 32'd115;
     memory[4940] = 32'd115;
     memory[4941] = 32'd179;
     memory[4942] = 32'd129;
     memory[4943] = 32'd4;
     memory[4944] = 32'd162;
     memory[4945] = 32'd233;
     memory[4946] = 32'd96;
     memory[4947] = 32'd148;
     memory[4948] = 32'd169;
     memory[4949] = 32'd77;
     memory[4950] = 32'd115;
     memory[4951] = 32'd141;
     memory[4952] = 32'd107;
     memory[4953] = 32'd71;
     memory[4954] = 32'd252;
     memory[4955] = 32'd182;
     memory[4956] = 32'd67;
     memory[4957] = 32'd36;
     memory[4958] = 32'd97;
     memory[4959] = 32'd25;
     memory[4960] = 32'd230;
     memory[4961] = 32'd55;
     memory[4962] = 32'd142;
     memory[4963] = 32'd194;
     memory[4964] = 32'd95;
     memory[4965] = 32'd121;
     memory[4966] = 32'd165;
     memory[4967] = 32'd230;
     memory[4968] = 32'd77;
     memory[4969] = 32'd226;
     memory[4970] = 32'd162;
     memory[4971] = 32'd237;
     memory[4972] = 32'd173;
     memory[4973] = 32'd230;
     memory[4974] = 32'd202;
     memory[4975] = 32'd102;
     memory[4976] = 32'd234;
     memory[4977] = 32'd99;
     memory[4978] = 32'd251;
     memory[4979] = 32'd152;
     memory[4980] = 32'd136;
     memory[4981] = 32'd32;
     memory[4982] = 32'd0;
     memory[4983] = 32'd210;
     memory[4984] = 32'd109;
     memory[4985] = 32'd55;
     memory[4986] = 32'd63;
     memory[4987] = 32'd173;
     memory[4988] = 32'd126;
     memory[4989] = 32'd165;
     memory[4990] = 32'd159;
     memory[4991] = 32'd85;
     memory[4992] = 32'd199;
     memory[4993] = 32'd57;
     memory[4994] = 32'd130;
     memory[4995] = 32'd193;
     memory[4996] = 32'd160;
     memory[4997] = 32'd24;
     memory[4998] = 32'd99;
     memory[4999] = 32'd252;
     memory[5000] = 32'd102;
     memory[5001] = 32'd58;
     memory[5002] = 32'd145;
     memory[5003] = 32'd18;
     memory[5004] = 32'd17;
     memory[5005] = 32'd116;
     memory[5006] = 32'd35;
     memory[5007] = 32'd107;
     memory[5008] = 32'd94;
     memory[5009] = 32'd211;
     memory[5010] = 32'd3;
     memory[5011] = 32'd75;
     memory[5012] = 32'd195;
     memory[5013] = 32'd181;
     memory[5014] = 32'd223;
     memory[5015] = 32'd186;
     memory[5016] = 32'd12;
     memory[5017] = 32'd238;
     memory[5018] = 32'd36;
     memory[5019] = 32'd107;
     memory[5020] = 32'd38;
     memory[5021] = 32'd46;
     memory[5022] = 32'd101;
     memory[5023] = 32'd233;
     memory[5024] = 32'd166;
     memory[5025] = 32'd130;
     memory[5026] = 32'd116;
     memory[5027] = 32'd179;
     memory[5028] = 32'd196;
     memory[5029] = 32'd13;
     memory[5030] = 32'd69;
     memory[5031] = 32'd82;
     memory[5032] = 32'd230;
     memory[5033] = 32'd175;
     memory[5034] = 32'd122;
     memory[5035] = 32'd26;
     memory[5036] = 32'd242;
     memory[5037] = 32'd231;
     memory[5038] = 32'd235;
     memory[5039] = 32'd218;
     memory[5040] = 32'd156;
     memory[5041] = 32'd57;
     memory[5042] = 32'd67;
     memory[5043] = 32'd160;
     memory[5044] = 32'd16;
     memory[5045] = 32'd186;
     memory[5046] = 32'd17;
     memory[5047] = 32'd197;
     memory[5048] = 32'd31;
     memory[5049] = 32'd167;
     memory[5050] = 32'd155;
     memory[5051] = 32'd26;
     memory[5052] = 32'd33;
     memory[5053] = 32'd89;
     memory[5054] = 32'd53;
     memory[5055] = 32'd69;
     memory[5056] = 32'd234;
     memory[5057] = 32'd234;
     memory[5058] = 32'd98;
     memory[5059] = 32'd203;
     memory[5060] = 32'd72;
     memory[5061] = 32'd129;
     memory[5062] = 32'd231;
     memory[5063] = 32'd91;
     memory[5064] = 32'd133;
     memory[5065] = 32'd89;
     memory[5066] = 32'd102;
     memory[5067] = 32'd149;
     memory[5068] = 32'd65;
     memory[5069] = 32'd233;
     memory[5070] = 32'd54;
     memory[5071] = 32'd29;
     memory[5072] = 32'd162;
     memory[5073] = 32'd251;
     memory[5074] = 32'd129;
     memory[5075] = 32'd143;
     memory[5076] = 32'd229;
     memory[5077] = 32'd127;
     memory[5078] = 32'd46;
     memory[5079] = 32'd140;
     memory[5080] = 32'd194;
     memory[5081] = 32'd173;
     memory[5082] = 32'd228;
     memory[5083] = 32'd129;
     memory[5084] = 32'd149;
     memory[5085] = 32'd104;
     memory[5086] = 32'd63;
     memory[5087] = 32'd237;
     memory[5088] = 32'd196;
     memory[5089] = 32'd68;
     memory[5090] = 32'd167;
     memory[5091] = 32'd55;
     memory[5092] = 32'd157;
     memory[5093] = 32'd138;
     memory[5094] = 32'd45;
     memory[5095] = 32'd174;
     memory[5096] = 32'd48;
     memory[5097] = 32'd242;
     memory[5098] = 32'd197;
     memory[5099] = 32'd126;
     memory[5100] = 32'd47;
     memory[5101] = 32'd173;
     memory[5102] = 32'd129;
     memory[5103] = 32'd198;
     memory[5104] = 32'd203;
     memory[5105] = 32'd204;
     memory[5106] = 32'd91;
     memory[5107] = 32'd250;
     memory[5108] = 32'd218;
     memory[5109] = 32'd200;
     memory[5110] = 32'd209;
     memory[5111] = 32'd121;
     memory[5112] = 32'd224;
     memory[5113] = 32'd133;
     memory[5114] = 32'd222;
     memory[5115] = 32'd223;
     memory[5116] = 32'd198;
     memory[5117] = 32'd84;
     memory[5118] = 32'd37;
     memory[5119] = 32'd5;
     memory[5120] = 32'd89;
     memory[5121] = 32'd84;
     memory[5122] = 32'd167;
     memory[5123] = 32'd26;
     memory[5124] = 32'd224;
     memory[5125] = 32'd3;
     memory[5126] = 32'd102;
     memory[5127] = 32'd210;
     memory[5128] = 32'd178;
     memory[5129] = 32'd1;
     memory[5130] = 32'd215;
     memory[5131] = 32'd166;
     memory[5132] = 32'd99;
     memory[5133] = 32'd51;
     memory[5134] = 32'd202;
     memory[5135] = 32'd181;
     memory[5136] = 32'd83;
     memory[5137] = 32'd57;
     memory[5138] = 32'd45;
     memory[5139] = 32'd252;
     memory[5140] = 32'd79;
     memory[5141] = 32'd100;
     memory[5142] = 32'd6;
     memory[5143] = 32'd225;
     memory[5144] = 32'd173;
     memory[5145] = 32'd252;
     memory[5146] = 32'd72;
     memory[5147] = 32'd239;
     memory[5148] = 32'd13;
     memory[5149] = 32'd242;
     memory[5150] = 32'd0;
     memory[5151] = 32'd123;
     memory[5152] = 32'd21;
     memory[5153] = 32'd38;
     memory[5154] = 32'd156;
     memory[5155] = 32'd155;
     memory[5156] = 32'd210;
     memory[5157] = 32'd246;
     memory[5158] = 32'd27;
     memory[5159] = 32'd152;
     memory[5160] = 32'd99;
     memory[5161] = 32'd134;
     memory[5162] = 32'd8;
     memory[5163] = 32'd208;
     memory[5164] = 32'd25;
     memory[5165] = 32'd140;
     memory[5166] = 32'd135;
     memory[5167] = 32'd114;
     memory[5168] = 32'd130;
     memory[5169] = 32'd204;
     memory[5170] = 32'd118;
     memory[5171] = 32'd180;
     memory[5172] = 32'd197;
     memory[5173] = 32'd100;
     memory[5174] = 32'd87;
     memory[5175] = 32'd247;
     memory[5176] = 32'd146;
     memory[5177] = 32'd123;
     memory[5178] = 32'd80;
     memory[5179] = 32'd118;
     memory[5180] = 32'd125;
     memory[5181] = 32'd35;
     memory[5182] = 32'd92;
     memory[5183] = 32'd182;
     memory[5184] = 32'd172;
     memory[5185] = 32'd191;
     memory[5186] = 32'd114;
     memory[5187] = 32'd89;
     memory[5188] = 32'd7;
     memory[5189] = 32'd220;
     memory[5190] = 32'd205;
     memory[5191] = 32'd187;
     memory[5192] = 32'd105;
     memory[5193] = 32'd154;
     memory[5194] = 32'd205;
     memory[5195] = 32'd32;
     memory[5196] = 32'd244;
     memory[5197] = 32'd18;
     memory[5198] = 32'd203;
     memory[5199] = 32'd192;
     memory[5200] = 32'd238;
     memory[5201] = 32'd252;
     memory[5202] = 32'd150;
     memory[5203] = 32'd108;
     memory[5204] = 32'd47;
     memory[5205] = 32'd192;
     memory[5206] = 32'd223;
     memory[5207] = 32'd253;
     memory[5208] = 32'd62;
     memory[5209] = 32'd36;
     memory[5210] = 32'd209;
     memory[5211] = 32'd111;
     memory[5212] = 32'd82;
     memory[5213] = 32'd74;
     memory[5214] = 32'd127;
     memory[5215] = 32'd218;
     memory[5216] = 32'd250;
     memory[5217] = 32'd82;
     memory[5218] = 32'd49;
     memory[5219] = 32'd65;
     memory[5220] = 32'd104;
     memory[5221] = 32'd22;
     memory[5222] = 32'd19;
     memory[5223] = 32'd250;
     memory[5224] = 32'd24;
     memory[5225] = 32'd9;
     memory[5226] = 32'd27;
     memory[5227] = 32'd96;
     memory[5228] = 32'd172;
     memory[5229] = 32'd92;
     memory[5230] = 32'd209;
     memory[5231] = 32'd3;
     memory[5232] = 32'd202;
     memory[5233] = 32'd93;
     memory[5234] = 32'd41;
     memory[5235] = 32'd88;
     memory[5236] = 32'd117;
     memory[5237] = 32'd194;
     memory[5238] = 32'd233;
     memory[5239] = 32'd227;
     memory[5240] = 32'd126;
     memory[5241] = 32'd56;
     memory[5242] = 32'd116;
     memory[5243] = 32'd181;
     memory[5244] = 32'd101;
     memory[5245] = 32'd191;
     memory[5246] = 32'd86;
     memory[5247] = 32'd244;
     memory[5248] = 32'd4;
     memory[5249] = 32'd96;
     memory[5250] = 32'd223;
     memory[5251] = 32'd87;
     memory[5252] = 32'd202;
     memory[5253] = 32'd140;
     memory[5254] = 32'd88;
     memory[5255] = 32'd65;
     memory[5256] = 32'd234;
     memory[5257] = 32'd78;
     memory[5258] = 32'd97;
     memory[5259] = 32'd92;
     memory[5260] = 32'd153;
     memory[5261] = 32'd93;
     memory[5262] = 32'd20;
     memory[5263] = 32'd119;
     memory[5264] = 32'd92;
     memory[5265] = 32'd169;
     memory[5266] = 32'd196;
     memory[5267] = 32'd59;
     memory[5268] = 32'd107;
     memory[5269] = 32'd17;
     memory[5270] = 32'd167;
     memory[5271] = 32'd98;
     memory[5272] = 32'd11;
     memory[5273] = 32'd137;
     memory[5274] = 32'd83;
     memory[5275] = 32'd22;
     memory[5276] = 32'd130;
     memory[5277] = 32'd232;
     memory[5278] = 32'd61;
     memory[5279] = 32'd10;
     memory[5280] = 32'd103;
     memory[5281] = 32'd176;
     memory[5282] = 32'd214;
     memory[5283] = 32'd134;
     memory[5284] = 32'd71;
     memory[5285] = 32'd209;
     memory[5286] = 32'd232;
     memory[5287] = 32'd20;
     memory[5288] = 32'd233;
     memory[5289] = 32'd15;
     memory[5290] = 32'd218;
     memory[5291] = 32'd222;
     memory[5292] = 32'd47;
     memory[5293] = 32'd213;
     memory[5294] = 32'd0;
     memory[5295] = 32'd65;
     memory[5296] = 32'd146;
     memory[5297] = 32'd249;
     memory[5298] = 32'd63;
     memory[5299] = 32'd94;
     memory[5300] = 32'd207;
     memory[5301] = 32'd9;
     memory[5302] = 32'd200;
     memory[5303] = 32'd248;
     memory[5304] = 32'd67;
     memory[5305] = 32'd247;
     memory[5306] = 32'd2;
     memory[5307] = 32'd20;
     memory[5308] = 32'd219;
     memory[5309] = 32'd197;
     memory[5310] = 32'd138;
     memory[5311] = 32'd36;
     memory[5312] = 32'd20;
     memory[5313] = 32'd46;
     memory[5314] = 32'd36;
     memory[5315] = 32'd37;
     memory[5316] = 32'd243;
     memory[5317] = 32'd230;
     memory[5318] = 32'd228;
     memory[5319] = 32'd131;
     memory[5320] = 32'd210;
     memory[5321] = 32'd174;
     memory[5322] = 32'd122;
     memory[5323] = 32'd12;
     memory[5324] = 32'd70;
     memory[5325] = 32'd213;
     memory[5326] = 32'd204;
     memory[5327] = 32'd235;
     memory[5328] = 32'd185;
     memory[5329] = 32'd109;
     memory[5330] = 32'd199;
     memory[5331] = 32'd136;
     memory[5332] = 32'd81;
     memory[5333] = 32'd11;
     memory[5334] = 32'd62;
     memory[5335] = 32'd28;
     memory[5336] = 32'd221;
     memory[5337] = 32'd98;
     memory[5338] = 32'd231;
     memory[5339] = 32'd210;
     memory[5340] = 32'd147;
     memory[5341] = 32'd143;
     memory[5342] = 32'd144;
     memory[5343] = 32'd213;
     memory[5344] = 32'd102;
     memory[5345] = 32'd4;
     memory[5346] = 32'd44;
     memory[5347] = 32'd51;
     memory[5348] = 32'd196;
     memory[5349] = 32'd67;
     memory[5350] = 32'd129;
     memory[5351] = 32'd151;
     memory[5352] = 32'd73;
     memory[5353] = 32'd67;
     memory[5354] = 32'd157;
     memory[5355] = 32'd102;
     memory[5356] = 32'd50;
     memory[5357] = 32'd169;
     memory[5358] = 32'd43;
     memory[5359] = 32'd212;
     memory[5360] = 32'd159;
     memory[5361] = 32'd189;
     memory[5362] = 32'd15;
     memory[5363] = 32'd155;
     memory[5364] = 32'd29;
     memory[5365] = 32'd109;
     memory[5366] = 32'd17;
     memory[5367] = 32'd140;
     memory[5368] = 32'd85;
     memory[5369] = 32'd206;
     memory[5370] = 32'd216;
     memory[5371] = 32'd208;
     memory[5372] = 32'd26;
     memory[5373] = 32'd59;
     memory[5374] = 32'd118;
     memory[5375] = 32'd239;
     memory[5376] = 32'd153;
     memory[5377] = 32'd136;
     memory[5378] = 32'd82;
     memory[5379] = 32'd120;
     memory[5380] = 32'd193;
     memory[5381] = 32'd232;
     memory[5382] = 32'd116;
     memory[5383] = 32'd14;
     memory[5384] = 32'd146;
     memory[5385] = 32'd138;
     memory[5386] = 32'd205;
     memory[5387] = 32'd219;
     memory[5388] = 32'd24;
     memory[5389] = 32'd28;
     memory[5390] = 32'd54;
     memory[5391] = 32'd234;
     memory[5392] = 32'd137;
     memory[5393] = 32'd209;
     memory[5394] = 32'd230;
     memory[5395] = 32'd184;
     memory[5396] = 32'd219;
     memory[5397] = 32'd160;
     memory[5398] = 32'd229;
     memory[5399] = 32'd40;
     memory[5400] = 32'd158;
     memory[5401] = 32'd222;
     memory[5402] = 32'd34;
     memory[5403] = 32'd14;
     memory[5404] = 32'd106;
     memory[5405] = 32'd48;
     memory[5406] = 32'd21;
     memory[5407] = 32'd35;
     memory[5408] = 32'd214;
     memory[5409] = 32'd243;
     memory[5410] = 32'd129;
     memory[5411] = 32'd155;
     memory[5412] = 32'd102;
     memory[5413] = 32'd236;
     memory[5414] = 32'd63;
     memory[5415] = 32'd40;
     memory[5416] = 32'd149;
     memory[5417] = 32'd103;
     memory[5418] = 32'd28;
     memory[5419] = 32'd10;
     memory[5420] = 32'd106;
     memory[5421] = 32'd73;
     memory[5422] = 32'd119;
     memory[5423] = 32'd202;
     memory[5424] = 32'd116;
     memory[5425] = 32'd91;
     memory[5426] = 32'd176;
     memory[5427] = 32'd19;
     memory[5428] = 32'd13;
     memory[5429] = 32'd163;
     memory[5430] = 32'd64;
     memory[5431] = 32'd136;
     memory[5432] = 32'd12;
     memory[5433] = 32'd249;
     memory[5434] = 32'd125;
     memory[5435] = 32'd76;
     memory[5436] = 32'd230;
     memory[5437] = 32'd185;
     memory[5438] = 32'd34;
     memory[5439] = 32'd251;
     memory[5440] = 32'd132;
     memory[5441] = 32'd159;
     memory[5442] = 32'd235;
     memory[5443] = 32'd144;
     memory[5444] = 32'd19;
     memory[5445] = 32'd11;
     memory[5446] = 32'd64;
     memory[5447] = 32'd181;
     memory[5448] = 32'd180;
     memory[5449] = 32'd216;
     memory[5450] = 32'd129;
     memory[5451] = 32'd213;
     memory[5452] = 32'd42;
     memory[5453] = 32'd0;
     memory[5454] = 32'd162;
     memory[5455] = 32'd89;
     memory[5456] = 32'd53;
     memory[5457] = 32'd158;
     memory[5458] = 32'd140;
     memory[5459] = 32'd69;
     memory[5460] = 32'd106;
     memory[5461] = 32'd29;
     memory[5462] = 32'd30;
     memory[5463] = 32'd131;
     memory[5464] = 32'd28;
     memory[5465] = 32'd99;
     memory[5466] = 32'd189;
     memory[5467] = 32'd225;
     memory[5468] = 32'd185;
     memory[5469] = 32'd32;
     memory[5470] = 32'd186;
     memory[5471] = 32'd69;
     memory[5472] = 32'd75;
     memory[5473] = 32'd163;
     memory[5474] = 32'd87;
     memory[5475] = 32'd212;
     memory[5476] = 32'd23;
     memory[5477] = 32'd203;
     memory[5478] = 32'd75;
     memory[5479] = 32'd236;
     memory[5480] = 32'd234;
     memory[5481] = 32'd217;
     memory[5482] = 32'd218;
     memory[5483] = 32'd236;
     memory[5484] = 32'd187;
     memory[5485] = 32'd69;
     memory[5486] = 32'd1;
     memory[5487] = 32'd166;
     memory[5488] = 32'd139;
     memory[5489] = 32'd17;
     memory[5490] = 32'd231;
     memory[5491] = 32'd38;
     memory[5492] = 32'd93;
     memory[5493] = 32'd22;
     memory[5494] = 32'd212;
     memory[5495] = 32'd26;
     memory[5496] = 32'd77;
     memory[5497] = 32'd248;
     memory[5498] = 32'd239;
     memory[5499] = 32'd128;
     memory[5500] = 32'd202;
     memory[5501] = 32'd155;
     memory[5502] = 32'd131;
     memory[5503] = 32'd42;
     memory[5504] = 32'd139;
     memory[5505] = 32'd173;
     memory[5506] = 32'd129;
     memory[5507] = 32'd217;
     memory[5508] = 32'd176;
     memory[5509] = 32'd28;
     memory[5510] = 32'd159;
     memory[5511] = 32'd157;
     memory[5512] = 32'd14;
     memory[5513] = 32'd16;
     memory[5514] = 32'd72;
     memory[5515] = 32'd48;
     memory[5516] = 32'd224;
     memory[5517] = 32'd220;
     memory[5518] = 32'd143;
     memory[5519] = 32'd250;
     memory[5520] = 32'd34;
     memory[5521] = 32'd161;
     memory[5522] = 32'd63;
     memory[5523] = 32'd197;
     memory[5524] = 32'd13;
     memory[5525] = 32'd126;
     memory[5526] = 32'd49;
     memory[5527] = 32'd162;
     memory[5528] = 32'd134;
     memory[5529] = 32'd70;
     memory[5530] = 32'd31;
     memory[5531] = 32'd128;
     memory[5532] = 32'd157;
     memory[5533] = 32'd49;
     memory[5534] = 32'd64;
     memory[5535] = 32'd82;
     memory[5536] = 32'd174;
     memory[5537] = 32'd151;
     memory[5538] = 32'd214;
     memory[5539] = 32'd61;
     memory[5540] = 32'd192;
     memory[5541] = 32'd203;
     memory[5542] = 32'd139;
     memory[5543] = 32'd69;
     memory[5544] = 32'd30;
     memory[5545] = 32'd50;
     memory[5546] = 32'd73;
     memory[5547] = 32'd74;
     memory[5548] = 32'd187;
     memory[5549] = 32'd8;
     memory[5550] = 32'd87;
     memory[5551] = 32'd157;
     memory[5552] = 32'd185;
     memory[5553] = 32'd241;
     memory[5554] = 32'd148;
     memory[5555] = 32'd123;
     memory[5556] = 32'd55;
     memory[5557] = 32'd252;
     memory[5558] = 32'd52;
     memory[5559] = 32'd37;
     memory[5560] = 32'd203;
     memory[5561] = 32'd162;
     memory[5562] = 32'd45;
     memory[5563] = 32'd23;
     memory[5564] = 32'd226;
     memory[5565] = 32'd202;
     memory[5566] = 32'd26;
     memory[5567] = 32'd29;
     memory[5568] = 32'd237;
     memory[5569] = 32'd135;
     memory[5570] = 32'd42;
     memory[5571] = 32'd164;
     memory[5572] = 32'd128;
     memory[5573] = 32'd21;
     memory[5574] = 32'd151;
     memory[5575] = 32'd63;
     memory[5576] = 32'd228;
     memory[5577] = 32'd183;
     memory[5578] = 32'd165;
     memory[5579] = 32'd167;
     memory[5580] = 32'd4;
     memory[5581] = 32'd211;
     memory[5582] = 32'd245;
     memory[5583] = 32'd62;
     memory[5584] = 32'd54;
     memory[5585] = 32'd235;
     memory[5586] = 32'd223;
     memory[5587] = 32'd61;
     memory[5588] = 32'd61;
     memory[5589] = 32'd48;
     memory[5590] = 32'd170;
     memory[5591] = 32'd213;
     memory[5592] = 32'd28;
     memory[5593] = 32'd218;
     memory[5594] = 32'd181;
     memory[5595] = 32'd221;
     memory[5596] = 32'd161;
     memory[5597] = 32'd65;
     memory[5598] = 32'd135;
     memory[5599] = 32'd185;
     memory[5600] = 32'd236;
     memory[5601] = 32'd19;
     memory[5602] = 32'd12;
     memory[5603] = 32'd225;
     memory[5604] = 32'd113;
     memory[5605] = 32'd53;
     memory[5606] = 32'd226;
     memory[5607] = 32'd72;
     memory[5608] = 32'd69;
     memory[5609] = 32'd105;
     memory[5610] = 32'd173;
     memory[5611] = 32'd116;
     memory[5612] = 32'd191;
     memory[5613] = 32'd4;
     memory[5614] = 32'd160;
     memory[5615] = 32'd233;
     memory[5616] = 32'd163;
     memory[5617] = 32'd199;
     memory[5618] = 32'd230;
     memory[5619] = 32'd29;
     memory[5620] = 32'd83;
     memory[5621] = 32'd23;
     memory[5622] = 32'd127;
     memory[5623] = 32'd113;
     memory[5624] = 32'd70;
     memory[5625] = 32'd204;
     memory[5626] = 32'd82;
     memory[5627] = 32'd209;
     memory[5628] = 32'd9;
     memory[5629] = 32'd63;
     memory[5630] = 32'd211;
     memory[5631] = 32'd111;
     memory[5632] = 32'd46;
     memory[5633] = 32'd160;
     memory[5634] = 32'd2;
     memory[5635] = 32'd171;
     memory[5636] = 32'd234;
     memory[5637] = 32'd102;
     memory[5638] = 32'd233;
     memory[5639] = 32'd52;
     memory[5640] = 32'd159;
     memory[5641] = 32'd137;
     memory[5642] = 32'd206;
     memory[5643] = 32'd77;
     memory[5644] = 32'd145;
     memory[5645] = 32'd236;
     memory[5646] = 32'd216;
     memory[5647] = 32'd55;
     memory[5648] = 32'd178;
     memory[5649] = 32'd182;
     memory[5650] = 32'd238;
     memory[5651] = 32'd222;
     memory[5652] = 32'd37;
     memory[5653] = 32'd120;
     memory[5654] = 32'd246;
     memory[5655] = 32'd180;
     memory[5656] = 32'd252;
     memory[5657] = 32'd12;
     memory[5658] = 32'd78;
     memory[5659] = 32'd232;
     memory[5660] = 32'd241;
     memory[5661] = 32'd116;
     memory[5662] = 32'd225;
     memory[5663] = 32'd163;
     memory[5664] = 32'd209;
     memory[5665] = 32'd49;
     memory[5666] = 32'd167;
     memory[5667] = 32'd159;
     memory[5668] = 32'd195;
     memory[5669] = 32'd238;
     memory[5670] = 32'd65;
     memory[5671] = 32'd245;
     memory[5672] = 32'd245;
     memory[5673] = 32'd85;
     memory[5674] = 32'd127;
     memory[5675] = 32'd55;
     memory[5676] = 32'd171;
     memory[5677] = 32'd80;
     memory[5678] = 32'd9;
     memory[5679] = 32'd95;
     memory[5680] = 32'd133;
     memory[5681] = 32'd58;
     memory[5682] = 32'd23;
     memory[5683] = 32'd69;
     memory[5684] = 32'd218;
     memory[5685] = 32'd203;
     memory[5686] = 32'd76;
     memory[5687] = 32'd163;
     memory[5688] = 32'd85;
     memory[5689] = 32'd137;
     memory[5690] = 32'd81;
     memory[5691] = 32'd124;
     memory[5692] = 32'd56;
     memory[5693] = 32'd151;
     memory[5694] = 32'd26;
     memory[5695] = 32'd102;
     memory[5696] = 32'd212;
     memory[5697] = 32'd74;
     memory[5698] = 32'd121;
     memory[5699] = 32'd13;
     memory[5700] = 32'd216;
     memory[5701] = 32'd64;
     memory[5702] = 32'd161;
     memory[5703] = 32'd207;
     memory[5704] = 32'd136;
     memory[5705] = 32'd6;
     memory[5706] = 32'd30;
     memory[5707] = 32'd79;
     memory[5708] = 32'd169;
     memory[5709] = 32'd66;
     memory[5710] = 32'd97;
     memory[5711] = 32'd76;
     memory[5712] = 32'd186;
     memory[5713] = 32'd202;
     memory[5714] = 32'd91;
     memory[5715] = 32'd19;
     memory[5716] = 32'd233;
     memory[5717] = 32'd161;
     memory[5718] = 32'd207;
     memory[5719] = 32'd24;
     memory[5720] = 32'd52;
     memory[5721] = 32'd151;
     memory[5722] = 32'd18;
     memory[5723] = 32'd174;
     memory[5724] = 32'd187;
     memory[5725] = 32'd235;
     memory[5726] = 32'd122;
     memory[5727] = 32'd86;
     memory[5728] = 32'd34;
     memory[5729] = 32'd141;
     memory[5730] = 32'd247;
     memory[5731] = 32'd107;
     memory[5732] = 32'd133;
     memory[5733] = 32'd206;
     memory[5734] = 32'd28;
     memory[5735] = 32'd53;
     memory[5736] = 32'd177;
     memory[5737] = 32'd104;
     memory[5738] = 32'd53;
     memory[5739] = 32'd53;
     memory[5740] = 32'd192;
     memory[5741] = 32'd1;
     memory[5742] = 32'd229;
     memory[5743] = 32'd218;
     memory[5744] = 32'd122;
     memory[5745] = 32'd151;
     memory[5746] = 32'd122;
     memory[5747] = 32'd23;
     memory[5748] = 32'd67;
     memory[5749] = 32'd204;
     memory[5750] = 32'd120;
     memory[5751] = 32'd0;
     memory[5752] = 32'd234;
     memory[5753] = 32'd5;
     memory[5754] = 32'd203;
     memory[5755] = 32'd213;
     memory[5756] = 32'd33;
     memory[5757] = 32'd135;
     memory[5758] = 32'd239;
     memory[5759] = 32'd44;
     memory[5760] = 32'd203;
     memory[5761] = 32'd127;
     memory[5762] = 32'd249;
     memory[5763] = 32'd26;
     memory[5764] = 32'd56;
     memory[5765] = 32'd45;
     memory[5766] = 32'd218;
     memory[5767] = 32'd111;
     memory[5768] = 32'd104;
     memory[5769] = 32'd252;
     memory[5770] = 32'd182;
     memory[5771] = 32'd148;
     memory[5772] = 32'd139;
     memory[5773] = 32'd0;
     memory[5774] = 32'd91;
     memory[5775] = 32'd172;
     memory[5776] = 32'd104;
     memory[5777] = 32'd138;
     memory[5778] = 32'd107;
     memory[5779] = 32'd216;
     memory[5780] = 32'd109;
     memory[5781] = 32'd165;
     memory[5782] = 32'd225;
     memory[5783] = 32'd89;
     memory[5784] = 32'd97;
     memory[5785] = 32'd108;
     memory[5786] = 32'd150;
     memory[5787] = 32'd54;
     memory[5788] = 32'd13;
     memory[5789] = 32'd178;
     memory[5790] = 32'd178;
     memory[5791] = 32'd204;
     memory[5792] = 32'd253;
     memory[5793] = 32'd52;
     memory[5794] = 32'd83;
     memory[5795] = 32'd65;
     memory[5796] = 32'd138;
     memory[5797] = 32'd55;
     memory[5798] = 32'd246;
     memory[5799] = 32'd82;
     memory[5800] = 32'd86;
     memory[5801] = 32'd212;
     memory[5802] = 32'd124;
     memory[5803] = 32'd227;
     memory[5804] = 32'd187;
     memory[5805] = 32'd197;
     memory[5806] = 32'd144;
     memory[5807] = 32'd201;
     memory[5808] = 32'd83;
     memory[5809] = 32'd74;
     memory[5810] = 32'd131;
     memory[5811] = 32'd135;
     memory[5812] = 32'd59;
     memory[5813] = 32'd204;
     memory[5814] = 32'd160;
     memory[5815] = 32'd210;
     memory[5816] = 32'd251;
     memory[5817] = 32'd156;
     memory[5818] = 32'd134;
     memory[5819] = 32'd69;
     memory[5820] = 32'd93;
     memory[5821] = 32'd231;
     memory[5822] = 32'd12;
     memory[5823] = 32'd97;
     memory[5824] = 32'd25;
     memory[5825] = 32'd110;
     memory[5826] = 32'd163;
     memory[5827] = 32'd112;
     memory[5828] = 32'd127;
     memory[5829] = 32'd55;
     memory[5830] = 32'd184;
     memory[5831] = 32'd145;
     memory[5832] = 32'd203;
     memory[5833] = 32'd166;
     memory[5834] = 32'd7;
     memory[5835] = 32'd110;
     memory[5836] = 32'd88;
     memory[5837] = 32'd116;
     memory[5838] = 32'd47;
     memory[5839] = 32'd57;
     memory[5840] = 32'd154;
     memory[5841] = 32'd58;
     memory[5842] = 32'd68;
     memory[5843] = 32'd192;
     memory[5844] = 32'd219;
     memory[5845] = 32'd124;
     memory[5846] = 32'd33;
     memory[5847] = 32'd90;
     memory[5848] = 32'd229;
     memory[5849] = 32'd241;
     memory[5850] = 32'd22;
     memory[5851] = 32'd204;
     memory[5852] = 32'd80;
     memory[5853] = 32'd193;
     memory[5854] = 32'd117;
     memory[5855] = 32'd177;
     memory[5856] = 32'd8;
     memory[5857] = 32'd51;
     memory[5858] = 32'd40;
     memory[5859] = 32'd45;
     memory[5860] = 32'd154;
     memory[5861] = 32'd4;
     memory[5862] = 32'd233;
     memory[5863] = 32'd162;
     memory[5864] = 32'd148;
     memory[5865] = 32'd231;
     memory[5866] = 32'd96;
     memory[5867] = 32'd218;
     memory[5868] = 32'd100;
     memory[5869] = 32'd244;
     memory[5870] = 32'd238;
     memory[5871] = 32'd16;
     memory[5872] = 32'd253;
     memory[5873] = 32'd76;
     memory[5874] = 32'd213;
     memory[5875] = 32'd254;
     memory[5876] = 32'd122;
     memory[5877] = 32'd91;
     memory[5878] = 32'd60;
     memory[5879] = 32'd158;
     memory[5880] = 32'd64;
     memory[5881] = 32'd101;
     memory[5882] = 32'd180;
     memory[5883] = 32'd46;
     memory[5884] = 32'd164;
     memory[5885] = 32'd57;
     memory[5886] = 32'd206;
     memory[5887] = 32'd158;
     memory[5888] = 32'd196;
     memory[5889] = 32'd80;
     memory[5890] = 32'd150;
     memory[5891] = 32'd20;
     memory[5892] = 32'd106;
     memory[5893] = 32'd92;
     memory[5894] = 32'd123;
     memory[5895] = 32'd122;
     memory[5896] = 32'd92;
     memory[5897] = 32'd157;
     memory[5898] = 32'd236;
     memory[5899] = 32'd79;
     memory[5900] = 32'd200;
     memory[5901] = 32'd103;
     memory[5902] = 32'd154;
     memory[5903] = 32'd201;
     memory[5904] = 32'd143;
     memory[5905] = 32'd93;
     memory[5906] = 32'd77;
     memory[5907] = 32'd144;
     memory[5908] = 32'd177;
     memory[5909] = 32'd207;
     memory[5910] = 32'd215;
     memory[5911] = 32'd57;
     memory[5912] = 32'd63;
     memory[5913] = 32'd48;
     memory[5914] = 32'd48;
     memory[5915] = 32'd145;
     memory[5916] = 32'd229;
     memory[5917] = 32'd86;
     memory[5918] = 32'd64;
     memory[5919] = 32'd109;
     memory[5920] = 32'd46;
     memory[5921] = 32'd41;
     memory[5922] = 32'd0;
     memory[5923] = 32'd44;
     memory[5924] = 32'd46;
     memory[5925] = 32'd5;
     memory[5926] = 32'd55;
     memory[5927] = 32'd178;
     memory[5928] = 32'd13;
     memory[5929] = 32'd24;
     memory[5930] = 32'd40;
     memory[5931] = 32'd69;
     memory[5932] = 32'd54;
     memory[5933] = 32'd96;
     memory[5934] = 32'd25;
     memory[5935] = 32'd81;
     memory[5936] = 32'd226;
     memory[5937] = 32'd71;
     memory[5938] = 32'd91;
     memory[5939] = 32'd122;
     memory[5940] = 32'd77;
     memory[5941] = 32'd126;
     memory[5942] = 32'd144;
     memory[5943] = 32'd221;
     memory[5944] = 32'd29;
     memory[5945] = 32'd212;
     memory[5946] = 32'd250;
     memory[5947] = 32'd108;
     memory[5948] = 32'd115;
     memory[5949] = 32'd211;
     memory[5950] = 32'd37;
     memory[5951] = 32'd185;
     memory[5952] = 32'd175;
     memory[5953] = 32'd59;
     memory[5954] = 32'd49;
     memory[5955] = 32'd126;
     memory[5956] = 32'd67;
     memory[5957] = 32'd29;
     memory[5958] = 32'd168;
     memory[5959] = 32'd112;
     memory[5960] = 32'd207;
     memory[5961] = 32'd168;
     memory[5962] = 32'd190;
     memory[5963] = 32'd127;
     memory[5964] = 32'd90;
     memory[5965] = 32'd195;
     memory[5966] = 32'd25;
     memory[5967] = 32'd40;
     memory[5968] = 32'd117;
     memory[5969] = 32'd31;
     memory[5970] = 32'd250;
     memory[5971] = 32'd244;
     memory[5972] = 32'd29;
     memory[5973] = 32'd251;
     memory[5974] = 32'd243;
     memory[5975] = 32'd153;
     memory[5976] = 32'd66;
     memory[5977] = 32'd168;
     memory[5978] = 32'd129;
     memory[5979] = 32'd144;
     memory[5980] = 32'd197;
     memory[5981] = 32'd0;
     memory[5982] = 32'd206;
     memory[5983] = 32'd73;
     memory[5984] = 32'd137;
     memory[5985] = 32'd252;
     memory[5986] = 32'd165;
     memory[5987] = 32'd173;
     memory[5988] = 32'd159;
     memory[5989] = 32'd244;
     memory[5990] = 32'd200;
     memory[5991] = 32'd234;
     memory[5992] = 32'd133;
     memory[5993] = 32'd205;
     memory[5994] = 32'd8;
     memory[5995] = 32'd224;
     memory[5996] = 32'd145;
     memory[5997] = 32'd28;
     memory[5998] = 32'd114;
     memory[5999] = 32'd158;
     memory[6000] = 32'd54;
     memory[6001] = 32'd187;
     memory[6002] = 32'd238;
     memory[6003] = 32'd252;
     memory[6004] = 32'd9;
     memory[6005] = 32'd212;
     memory[6006] = 32'd145;
     memory[6007] = 32'd244;
     memory[6008] = 32'd2;
     memory[6009] = 32'd149;
     memory[6010] = 32'd83;
     memory[6011] = 32'd150;
     memory[6012] = 32'd71;
     memory[6013] = 32'd98;
     memory[6014] = 32'd24;
     memory[6015] = 32'd85;
     memory[6016] = 32'd122;
     memory[6017] = 32'd233;
     memory[6018] = 32'd214;
     memory[6019] = 32'd15;
     memory[6020] = 32'd109;
     memory[6021] = 32'd60;
     memory[6022] = 32'd170;
     memory[6023] = 32'd238;
     memory[6024] = 32'd72;
     memory[6025] = 32'd44;
     memory[6026] = 32'd190;
     memory[6027] = 32'd34;
     memory[6028] = 32'd76;
     memory[6029] = 32'd166;
     memory[6030] = 32'd177;
     memory[6031] = 32'd115;
     memory[6032] = 32'd57;
     memory[6033] = 32'd209;
     memory[6034] = 32'd96;
     memory[6035] = 32'd241;
     memory[6036] = 32'd5;
     memory[6037] = 32'd130;
     memory[6038] = 32'd149;
     memory[6039] = 32'd64;
     memory[6040] = 32'd233;
     memory[6041] = 32'd27;
     memory[6042] = 32'd63;
     memory[6043] = 32'd189;
     memory[6044] = 32'd96;
     memory[6045] = 32'd177;
     memory[6046] = 32'd152;
     memory[6047] = 32'd85;
     memory[6048] = 32'd223;
     memory[6049] = 32'd217;
     memory[6050] = 32'd59;
     memory[6051] = 32'd222;
     memory[6052] = 32'd155;
     memory[6053] = 32'd2;
     memory[6054] = 32'd131;
     memory[6055] = 32'd162;
     memory[6056] = 32'd19;
     memory[6057] = 32'd26;
     memory[6058] = 32'd95;
     memory[6059] = 32'd170;
     memory[6060] = 32'd226;
     memory[6061] = 32'd188;
     memory[6062] = 32'd138;
     memory[6063] = 32'd103;
     memory[6064] = 32'd146;
     memory[6065] = 32'd154;
     memory[6066] = 32'd150;
     memory[6067] = 32'd156;
     memory[6068] = 32'd52;
     memory[6069] = 32'd150;
     memory[6070] = 32'd165;
     memory[6071] = 32'd119;
     memory[6072] = 32'd15;
     memory[6073] = 32'd148;
     memory[6074] = 32'd65;
     memory[6075] = 32'd152;
     memory[6076] = 32'd142;
     memory[6077] = 32'd15;
     memory[6078] = 32'd84;
     memory[6079] = 32'd109;
     memory[6080] = 32'd252;
     memory[6081] = 32'd197;
     memory[6082] = 32'd225;
     memory[6083] = 32'd65;
     memory[6084] = 32'd64;
     memory[6085] = 32'd64;
     memory[6086] = 32'd110;
     memory[6087] = 32'd6;
     memory[6088] = 32'd45;
     memory[6089] = 32'd160;
     memory[6090] = 32'd111;
     memory[6091] = 32'd67;
     memory[6092] = 32'd52;
     memory[6093] = 32'd22;
     memory[6094] = 32'd11;
     memory[6095] = 32'd152;
     memory[6096] = 32'd6;
     memory[6097] = 32'd213;
     memory[6098] = 32'd59;
     memory[6099] = 32'd66;
     memory[6100] = 32'd92;
     memory[6101] = 32'd31;
     memory[6102] = 32'd235;
     memory[6103] = 32'd24;
     memory[6104] = 32'd102;
     memory[6105] = 32'd99;
     memory[6106] = 32'd216;
     memory[6107] = 32'd92;
     memory[6108] = 32'd87;
     memory[6109] = 32'd231;
     memory[6110] = 32'd170;
     memory[6111] = 32'd153;
     memory[6112] = 32'd192;
     memory[6113] = 32'd50;
     memory[6114] = 32'd204;
     memory[6115] = 32'd92;
     memory[6116] = 32'd165;
     memory[6117] = 32'd139;
     memory[6118] = 32'd1;
     memory[6119] = 32'd214;
     memory[6120] = 32'd196;
     memory[6121] = 32'd57;
     memory[6122] = 32'd129;
     memory[6123] = 32'd98;
     memory[6124] = 32'd87;
     memory[6125] = 32'd208;
     memory[6126] = 32'd125;
     memory[6127] = 32'd91;
     memory[6128] = 32'd245;
     memory[6129] = 32'd115;
     memory[6130] = 32'd168;
     memory[6131] = 32'd72;
     memory[6132] = 32'd43;
     memory[6133] = 32'd159;
     memory[6134] = 32'd198;
     memory[6135] = 32'd190;
     memory[6136] = 32'd196;
     memory[6137] = 32'd163;
     memory[6138] = 32'd66;
     memory[6139] = 32'd164;
     memory[6140] = 32'd25;
     memory[6141] = 32'd223;
     memory[6142] = 32'd10;
     memory[6143] = 32'd163;
     memory[6144] = 32'd1;
     memory[6145] = 32'd71;
     memory[6146] = 32'd180;
     memory[6147] = 32'd8;
     memory[6148] = 32'd27;
     memory[6149] = 32'd133;
     memory[6150] = 32'd34;
     memory[6151] = 32'd195;
     memory[6152] = 32'd206;
     memory[6153] = 32'd42;
     memory[6154] = 32'd154;
     memory[6155] = 32'd81;
     memory[6156] = 32'd31;
     memory[6157] = 32'd105;
     memory[6158] = 32'd236;
     memory[6159] = 32'd59;
     memory[6160] = 32'd83;
     memory[6161] = 32'd99;
     memory[6162] = 32'd38;
     memory[6163] = 32'd254;
     memory[6164] = 32'd170;
     memory[6165] = 32'd41;
     memory[6166] = 32'd47;
     memory[6167] = 32'd236;
     memory[6168] = 32'd231;
     memory[6169] = 32'd32;
     memory[6170] = 32'd166;
     memory[6171] = 32'd60;
     memory[6172] = 32'd213;
     memory[6173] = 32'd27;
     memory[6174] = 32'd120;
     memory[6175] = 32'd166;
     memory[6176] = 32'd247;
     memory[6177] = 32'd213;
     memory[6178] = 32'd242;
     memory[6179] = 32'd227;
     memory[6180] = 32'd98;
     memory[6181] = 32'd132;
     memory[6182] = 32'd92;
     memory[6183] = 32'd48;
     memory[6184] = 32'd110;
     memory[6185] = 32'd185;
     memory[6186] = 32'd183;
     memory[6187] = 32'd226;
     memory[6188] = 32'd60;
     memory[6189] = 32'd134;
     memory[6190] = 32'd251;
     memory[6191] = 32'd127;
     memory[6192] = 32'd33;
     memory[6193] = 32'd87;
     memory[6194] = 32'd105;
     memory[6195] = 32'd110;
     memory[6196] = 32'd220;
     memory[6197] = 32'd27;
     memory[6198] = 32'd76;
     memory[6199] = 32'd132;
     memory[6200] = 32'd150;
     memory[6201] = 32'd105;
     memory[6202] = 32'd100;
     memory[6203] = 32'd17;
     memory[6204] = 32'd98;
     memory[6205] = 32'd183;
     memory[6206] = 32'd35;
     memory[6207] = 32'd254;
     memory[6208] = 32'd4;
     memory[6209] = 32'd234;
     memory[6210] = 32'd154;
     memory[6211] = 32'd25;
     memory[6212] = 32'd113;
     memory[6213] = 32'd231;
     memory[6214] = 32'd14;
     memory[6215] = 32'd251;
     memory[6216] = 32'd74;
     memory[6217] = 32'd2;
     memory[6218] = 32'd8;
     memory[6219] = 32'd63;
     memory[6220] = 32'd58;
     memory[6221] = 32'd73;
     memory[6222] = 32'd27;
     memory[6223] = 32'd52;
     memory[6224] = 32'd167;
     memory[6225] = 32'd78;
     memory[6226] = 32'd230;
     memory[6227] = 32'd171;
     memory[6228] = 32'd101;
     memory[6229] = 32'd172;
     memory[6230] = 32'd51;
     memory[6231] = 32'd10;
     memory[6232] = 32'd27;
     memory[6233] = 32'd119;
     memory[6234] = 32'd214;
     memory[6235] = 32'd49;
     memory[6236] = 32'd61;
     memory[6237] = 32'd36;
     memory[6238] = 32'd231;
     memory[6239] = 32'd94;
     memory[6240] = 32'd45;
     memory[6241] = 32'd170;
     memory[6242] = 32'd149;
     memory[6243] = 32'd250;
     memory[6244] = 32'd45;
     memory[6245] = 32'd118;
     memory[6246] = 32'd124;
     memory[6247] = 32'd69;
     memory[6248] = 32'd32;
     memory[6249] = 32'd22;
     memory[6250] = 32'd122;
     memory[6251] = 32'd172;
     memory[6252] = 32'd18;
     memory[6253] = 32'd10;
     memory[6254] = 32'd107;
     memory[6255] = 32'd164;
     memory[6256] = 32'd113;
     memory[6257] = 32'd139;
     memory[6258] = 32'd130;
     memory[6259] = 32'd212;
     memory[6260] = 32'd72;
     memory[6261] = 32'd117;
     memory[6262] = 32'd102;
     memory[6263] = 32'd88;
     memory[6264] = 32'd169;
     memory[6265] = 32'd252;
     memory[6266] = 32'd122;
     memory[6267] = 32'd182;
     memory[6268] = 32'd126;
     memory[6269] = 32'd106;
     memory[6270] = 32'd77;
     memory[6271] = 32'd160;
     memory[6272] = 32'd156;
     memory[6273] = 32'd143;
     memory[6274] = 32'd120;
     memory[6275] = 32'd130;
     memory[6276] = 32'd91;
     memory[6277] = 32'd218;
     memory[6278] = 32'd147;
     memory[6279] = 32'd123;
     memory[6280] = 32'd30;
     memory[6281] = 32'd121;
     memory[6282] = 32'd70;
     memory[6283] = 32'd194;
     memory[6284] = 32'd136;
     memory[6285] = 32'd194;
     memory[6286] = 32'd29;
     memory[6287] = 32'd53;
     memory[6288] = 32'd12;
     memory[6289] = 32'd127;
     memory[6290] = 32'd142;
     memory[6291] = 32'd112;
     memory[6292] = 32'd75;
     memory[6293] = 32'd139;
     memory[6294] = 32'd93;
     memory[6295] = 32'd229;
     memory[6296] = 32'd182;
     memory[6297] = 32'd158;
     memory[6298] = 32'd22;
     memory[6299] = 32'd25;
     memory[6300] = 32'd118;
     memory[6301] = 32'd102;
     memory[6302] = 32'd186;
     memory[6303] = 32'd185;
     memory[6304] = 32'd204;
     memory[6305] = 32'd116;
     memory[6306] = 32'd89;
     memory[6307] = 32'd12;
     memory[6308] = 32'd167;
     memory[6309] = 32'd153;
     memory[6310] = 32'd161;
     memory[6311] = 32'd18;
     memory[6312] = 32'd125;
     memory[6313] = 32'd126;
     memory[6314] = 32'd213;
     memory[6315] = 32'd8;
     memory[6316] = 32'd110;
     memory[6317] = 32'd130;
     memory[6318] = 32'd168;
     memory[6319] = 32'd176;
     memory[6320] = 32'd169;
     memory[6321] = 32'd205;
     memory[6322] = 32'd16;
     memory[6323] = 32'd233;
     memory[6324] = 32'd66;
     memory[6325] = 32'd224;
     memory[6326] = 32'd128;
     memory[6327] = 32'd204;
     memory[6328] = 32'd42;
     memory[6329] = 32'd172;
     memory[6330] = 32'd119;
     memory[6331] = 32'd18;
     memory[6332] = 32'd11;
     memory[6333] = 32'd26;
     memory[6334] = 32'd12;
     memory[6335] = 32'd140;
     memory[6336] = 32'd163;
     memory[6337] = 32'd235;
     memory[6338] = 32'd89;
     memory[6339] = 32'd21;
     memory[6340] = 32'd252;
     memory[6341] = 32'd71;
     memory[6342] = 32'd195;
     memory[6343] = 32'd2;
     memory[6344] = 32'd224;
     memory[6345] = 32'd124;
     memory[6346] = 32'd7;
     memory[6347] = 32'd120;
     memory[6348] = 32'd60;
     memory[6349] = 32'd215;
     memory[6350] = 32'd30;
     memory[6351] = 32'd171;
     memory[6352] = 32'd71;
     memory[6353] = 32'd175;
     memory[6354] = 32'd96;
     memory[6355] = 32'd179;
     memory[6356] = 32'd146;
     memory[6357] = 32'd194;
     memory[6358] = 32'd143;
     memory[6359] = 32'd163;
     memory[6360] = 32'd28;
     memory[6361] = 32'd114;
     memory[6362] = 32'd252;
     memory[6363] = 32'd225;
     memory[6364] = 32'd230;
     memory[6365] = 32'd155;
     memory[6366] = 32'd95;
     memory[6367] = 32'd56;
     memory[6368] = 32'd198;
     memory[6369] = 32'd236;
     memory[6370] = 32'd210;
     memory[6371] = 32'd240;
     memory[6372] = 32'd112;
     memory[6373] = 32'd242;
     memory[6374] = 32'd210;
     memory[6375] = 32'd223;
     memory[6376] = 32'd219;
     memory[6377] = 32'd126;
     memory[6378] = 32'd249;
     memory[6379] = 32'd158;
     memory[6380] = 32'd73;
     memory[6381] = 32'd119;
     memory[6382] = 32'd84;
     memory[6383] = 32'd183;
     memory[6384] = 32'd0;
     memory[6385] = 32'd20;
     memory[6386] = 32'd194;
     memory[6387] = 32'd124;
     memory[6388] = 32'd88;
     memory[6389] = 32'd216;
     memory[6390] = 32'd165;
     memory[6391] = 32'd114;
     memory[6392] = 32'd69;
     memory[6393] = 32'd164;
     memory[6394] = 32'd124;
     memory[6395] = 32'd231;
     memory[6396] = 32'd50;
     memory[6397] = 32'd67;
     memory[6398] = 32'd156;
     memory[6399] = 32'd242;
     memory[6400] = 32'd152;
     memory[6401] = 32'd94;
     memory[6402] = 32'd198;
     memory[6403] = 32'd234;
     memory[6404] = 32'd50;
     memory[6405] = 32'd233;
     memory[6406] = 32'd216;
     memory[6407] = 32'd32;
     memory[6408] = 32'd235;
     memory[6409] = 32'd30;
     memory[6410] = 32'd108;
     memory[6411] = 32'd208;
     memory[6412] = 32'd228;
     memory[6413] = 32'd124;
     memory[6414] = 32'd87;
     memory[6415] = 32'd127;
     memory[6416] = 32'd192;
     memory[6417] = 32'd27;
     memory[6418] = 32'd58;
     memory[6419] = 32'd59;
     memory[6420] = 32'd126;
     memory[6421] = 32'd254;
     memory[6422] = 32'd92;
     memory[6423] = 32'd5;
     memory[6424] = 32'd67;
     memory[6425] = 32'd197;
     memory[6426] = 32'd165;
     memory[6427] = 32'd43;
     memory[6428] = 32'd7;
     memory[6429] = 32'd112;
     memory[6430] = 32'd129;
     memory[6431] = 32'd85;
     memory[6432] = 32'd206;
     memory[6433] = 32'd111;
     memory[6434] = 32'd25;
     memory[6435] = 32'd216;
     memory[6436] = 32'd51;
     memory[6437] = 32'd61;
     memory[6438] = 32'd131;
     memory[6439] = 32'd52;
     memory[6440] = 32'd200;
     memory[6441] = 32'd232;
     memory[6442] = 32'd16;
     memory[6443] = 32'd160;
     memory[6444] = 32'd166;
     memory[6445] = 32'd107;
     memory[6446] = 32'd178;
     memory[6447] = 32'd220;
     memory[6448] = 32'd114;
     memory[6449] = 32'd119;
     memory[6450] = 32'd149;
     memory[6451] = 32'd253;
     memory[6452] = 32'd81;
     memory[6453] = 32'd201;
     memory[6454] = 32'd209;
     memory[6455] = 32'd66;
     memory[6456] = 32'd155;
     memory[6457] = 32'd91;
     memory[6458] = 32'd198;
     memory[6459] = 32'd138;
     memory[6460] = 32'd83;
     memory[6461] = 32'd35;
     memory[6462] = 32'd138;
     memory[6463] = 32'd189;
     memory[6464] = 32'd180;
     memory[6465] = 32'd27;
     memory[6466] = 32'd158;
     memory[6467] = 32'd22;
     memory[6468] = 32'd251;
     memory[6469] = 32'd40;
     memory[6470] = 32'd161;
     memory[6471] = 32'd180;
     memory[6472] = 32'd135;
     memory[6473] = 32'd68;
     memory[6474] = 32'd126;
     memory[6475] = 32'd203;
     memory[6476] = 32'd60;
     memory[6477] = 32'd213;
     memory[6478] = 32'd185;
     memory[6479] = 32'd6;
     memory[6480] = 32'd136;
     memory[6481] = 32'd30;
     memory[6482] = 32'd100;
     memory[6483] = 32'd128;
     memory[6484] = 32'd7;
     memory[6485] = 32'd13;
     memory[6486] = 32'd18;
     memory[6487] = 32'd160;
     memory[6488] = 32'd197;
     memory[6489] = 32'd212;
     memory[6490] = 32'd244;
     memory[6491] = 32'd127;
     memory[6492] = 32'd173;
     memory[6493] = 32'd80;
     memory[6494] = 32'd134;
     memory[6495] = 32'd104;
     memory[6496] = 32'd101;
     memory[6497] = 32'd9;
     memory[6498] = 32'd15;
     memory[6499] = 32'd195;
     memory[6500] = 32'd223;
     memory[6501] = 32'd141;
     memory[6502] = 32'd134;
     memory[6503] = 32'd75;
     memory[6504] = 32'd112;
     memory[6505] = 32'd3;
     memory[6506] = 32'd92;
     memory[6507] = 32'd81;
     memory[6508] = 32'd2;
     memory[6509] = 32'd244;
     memory[6510] = 32'd16;
     memory[6511] = 32'd70;
     memory[6512] = 32'd164;
     memory[6513] = 32'd84;
     memory[6514] = 32'd93;
     memory[6515] = 32'd146;
     memory[6516] = 32'd146;
     memory[6517] = 32'd180;
     memory[6518] = 32'd241;
     memory[6519] = 32'd1;
     memory[6520] = 32'd226;
     memory[6521] = 32'd183;
     memory[6522] = 32'd43;
     memory[6523] = 32'd136;
     memory[6524] = 32'd143;
     memory[6525] = 32'd222;
     memory[6526] = 32'd143;
     memory[6527] = 32'd237;
     memory[6528] = 32'd169;
     memory[6529] = 32'd218;
     memory[6530] = 32'd5;
     memory[6531] = 32'd187;
     memory[6532] = 32'd42;
     memory[6533] = 32'd93;
     memory[6534] = 32'd215;
     memory[6535] = 32'd148;
     memory[6536] = 32'd54;
     memory[6537] = 32'd152;
     memory[6538] = 32'd228;
     memory[6539] = 32'd130;
     memory[6540] = 32'd3;
     memory[6541] = 32'd156;
     memory[6542] = 32'd172;
     memory[6543] = 32'd239;
     memory[6544] = 32'd42;
     memory[6545] = 32'd232;
     memory[6546] = 32'd233;
     memory[6547] = 32'd76;
     memory[6548] = 32'd88;
     memory[6549] = 32'd234;
     memory[6550] = 32'd64;
     memory[6551] = 32'd123;
     memory[6552] = 32'd169;
     memory[6553] = 32'd201;
     memory[6554] = 32'd165;
     memory[6555] = 32'd147;
     memory[6556] = 32'd73;
     memory[6557] = 32'd214;
     memory[6558] = 32'd97;
     memory[6559] = 32'd87;
     memory[6560] = 32'd43;
     memory[6561] = 32'd146;
     memory[6562] = 32'd88;
     memory[6563] = 32'd214;
     memory[6564] = 32'd98;
     memory[6565] = 32'd99;
     memory[6566] = 32'd156;
     memory[6567] = 32'd248;
     memory[6568] = 32'd132;
     memory[6569] = 32'd157;
     memory[6570] = 32'd215;
     memory[6571] = 32'd57;
     memory[6572] = 32'd2;
     memory[6573] = 32'd71;
     memory[6574] = 32'd0;
     memory[6575] = 32'd33;
     memory[6576] = 32'd126;
     memory[6577] = 32'd190;
     memory[6578] = 32'd234;
     memory[6579] = 32'd195;
     memory[6580] = 32'd28;
     memory[6581] = 32'd4;
     memory[6582] = 32'd36;
     memory[6583] = 32'd214;
     memory[6584] = 32'd88;
     memory[6585] = 32'd36;
     memory[6586] = 32'd205;
     memory[6587] = 32'd180;
     memory[6588] = 32'd47;
     memory[6589] = 32'd233;
     memory[6590] = 32'd232;
     memory[6591] = 32'd29;
     memory[6592] = 32'd109;
     memory[6593] = 32'd18;
     memory[6594] = 32'd136;
     memory[6595] = 32'd216;
     memory[6596] = 32'd106;
     memory[6597] = 32'd76;
     memory[6598] = 32'd188;
     memory[6599] = 32'd70;
     memory[6600] = 32'd207;
     memory[6601] = 32'd101;
     memory[6602] = 32'd21;
     memory[6603] = 32'd68;
     memory[6604] = 32'd34;
     memory[6605] = 32'd245;
     memory[6606] = 32'd233;
     memory[6607] = 32'd43;
     memory[6608] = 32'd137;
     memory[6609] = 32'd215;
     memory[6610] = 32'd236;
     memory[6611] = 32'd189;
     memory[6612] = 32'd0;
     memory[6613] = 32'd240;
     memory[6614] = 32'd217;
     memory[6615] = 32'd28;
     memory[6616] = 32'd72;
     memory[6617] = 32'd36;
     memory[6618] = 32'd47;
     memory[6619] = 32'd115;
     memory[6620] = 32'd88;
     memory[6621] = 32'd193;
     memory[6622] = 32'd152;
     memory[6623] = 32'd87;
     memory[6624] = 32'd174;
     memory[6625] = 32'd79;
     memory[6626] = 32'd117;
     memory[6627] = 32'd170;
     memory[6628] = 32'd79;
     memory[6629] = 32'd9;
     memory[6630] = 32'd83;
     memory[6631] = 32'd138;
     memory[6632] = 32'd108;
     memory[6633] = 32'd57;
     memory[6634] = 32'd195;
     memory[6635] = 32'd186;
     memory[6636] = 32'd211;
     memory[6637] = 32'd3;
     memory[6638] = 32'd251;
     memory[6639] = 32'd80;
     memory[6640] = 32'd157;
     memory[6641] = 32'd5;
     memory[6642] = 32'd33;
     memory[6643] = 32'd147;
     memory[6644] = 32'd135;
     memory[6645] = 32'd27;
     memory[6646] = 32'd83;
     memory[6647] = 32'd138;
     memory[6648] = 32'd99;
     memory[6649] = 32'd98;
     memory[6650] = 32'd124;
     memory[6651] = 32'd29;
     memory[6652] = 32'd10;
     memory[6653] = 32'd74;
     memory[6654] = 32'd194;
     memory[6655] = 32'd96;
     memory[6656] = 32'd146;
     memory[6657] = 32'd209;
     memory[6658] = 32'd131;
     memory[6659] = 32'd171;
     memory[6660] = 32'd181;
     memory[6661] = 32'd12;
     memory[6662] = 32'd57;
     memory[6663] = 32'd112;
     memory[6664] = 32'd180;
     memory[6665] = 32'd3;
     memory[6666] = 32'd135;
     memory[6667] = 32'd18;
     memory[6668] = 32'd91;
     memory[6669] = 32'd72;
     memory[6670] = 32'd217;
     memory[6671] = 32'd83;
     memory[6672] = 32'd18;
     memory[6673] = 32'd201;
     memory[6674] = 32'd212;
     memory[6675] = 32'd182;
     memory[6676] = 32'd52;
     memory[6677] = 32'd72;
     memory[6678] = 32'd134;
     memory[6679] = 32'd40;
     memory[6680] = 32'd95;
     memory[6681] = 32'd25;
     memory[6682] = 32'd90;
     memory[6683] = 32'd252;
     memory[6684] = 32'd192;
     memory[6685] = 32'd193;
     memory[6686] = 32'd75;
     memory[6687] = 32'd212;
     memory[6688] = 32'd6;
     memory[6689] = 32'd140;
     memory[6690] = 32'd114;
     memory[6691] = 32'd182;
     memory[6692] = 32'd53;
     memory[6693] = 32'd118;
     memory[6694] = 32'd127;
     memory[6695] = 32'd16;
     memory[6696] = 32'd78;
     memory[6697] = 32'd31;
     memory[6698] = 32'd75;
     memory[6699] = 32'd135;
     memory[6700] = 32'd221;
     memory[6701] = 32'd193;
     memory[6702] = 32'd204;
     memory[6703] = 32'd1;
     memory[6704] = 32'd134;
     memory[6705] = 32'd84;
     memory[6706] = 32'd183;
     memory[6707] = 32'd123;
     memory[6708] = 32'd27;
     memory[6709] = 32'd62;
     memory[6710] = 32'd97;
     memory[6711] = 32'd32;
     memory[6712] = 32'd164;
     memory[6713] = 32'd120;
     memory[6714] = 32'd99;
     memory[6715] = 32'd57;
     memory[6716] = 32'd123;
     memory[6717] = 32'd68;
     memory[6718] = 32'd222;
     memory[6719] = 32'd242;
     memory[6720] = 32'd154;
     memory[6721] = 32'd242;
     memory[6722] = 32'd4;
     memory[6723] = 32'd188;
     memory[6724] = 32'd249;
     memory[6725] = 32'd212;
     memory[6726] = 32'd158;
     memory[6727] = 32'd101;
     memory[6728] = 32'd5;
     memory[6729] = 32'd16;
     memory[6730] = 32'd4;
     memory[6731] = 32'd34;
     memory[6732] = 32'd95;
     memory[6733] = 32'd237;
     memory[6734] = 32'd8;
     memory[6735] = 32'd139;
     memory[6736] = 32'd4;
     memory[6737] = 32'd108;
     memory[6738] = 32'd124;
     memory[6739] = 32'd53;
     memory[6740] = 32'd10;
     memory[6741] = 32'd101;
     memory[6742] = 32'd51;
     memory[6743] = 32'd197;
     memory[6744] = 32'd124;
     memory[6745] = 32'd130;
     memory[6746] = 32'd152;
     memory[6747] = 32'd238;
     memory[6748] = 32'd101;
     memory[6749] = 32'd190;
     memory[6750] = 32'd248;
     memory[6751] = 32'd37;
     memory[6752] = 32'd37;
     memory[6753] = 32'd37;
     memory[6754] = 32'd205;
     memory[6755] = 32'd7;
     memory[6756] = 32'd117;
     memory[6757] = 32'd9;
     memory[6758] = 32'd111;
     memory[6759] = 32'd47;
     memory[6760] = 32'd163;
     memory[6761] = 32'd25;
     memory[6762] = 32'd59;
     memory[6763] = 32'd183;
     memory[6764] = 32'd24;
     memory[6765] = 32'd190;
     memory[6766] = 32'd172;
     memory[6767] = 32'd160;
     memory[6768] = 32'd38;
     memory[6769] = 32'd196;
     memory[6770] = 32'd5;
     memory[6771] = 32'd159;
     memory[6772] = 32'd109;
     memory[6773] = 32'd138;
     memory[6774] = 32'd209;
     memory[6775] = 32'd114;
     memory[6776] = 32'd140;
     memory[6777] = 32'd6;
     memory[6778] = 32'd60;
     memory[6779] = 32'd240;
     memory[6780] = 32'd174;
     memory[6781] = 32'd85;
     memory[6782] = 32'd175;
     memory[6783] = 32'd252;
     memory[6784] = 32'd165;
     memory[6785] = 32'd83;
     memory[6786] = 32'd100;
     memory[6787] = 32'd181;
     memory[6788] = 32'd56;
     memory[6789] = 32'd199;
     memory[6790] = 32'd205;
     memory[6791] = 32'd100;
     memory[6792] = 32'd220;
     memory[6793] = 32'd163;
     memory[6794] = 32'd243;
     memory[6795] = 32'd166;
     memory[6796] = 32'd224;
     memory[6797] = 32'd124;
     memory[6798] = 32'd103;
     memory[6799] = 32'd124;
     memory[6800] = 32'd164;
     memory[6801] = 32'd172;
     memory[6802] = 32'd245;
     memory[6803] = 32'd28;
     memory[6804] = 32'd10;
     memory[6805] = 32'd6;
     memory[6806] = 32'd135;
     memory[6807] = 32'd50;
     memory[6808] = 32'd140;
     memory[6809] = 32'd169;
     memory[6810] = 32'd82;
     memory[6811] = 32'd141;
     memory[6812] = 32'd85;
     memory[6813] = 32'd194;
     memory[6814] = 32'd144;
     memory[6815] = 32'd45;
     memory[6816] = 32'd35;
     memory[6817] = 32'd125;
     memory[6818] = 32'd249;
     memory[6819] = 32'd129;
     memory[6820] = 32'd169;
     memory[6821] = 32'd133;
     memory[6822] = 32'd22;
     memory[6823] = 32'd191;
     memory[6824] = 32'd105;
     memory[6825] = 32'd195;
     memory[6826] = 32'd78;
     memory[6827] = 32'd167;
     memory[6828] = 32'd103;
     memory[6829] = 32'd153;
     memory[6830] = 32'd58;
     memory[6831] = 32'd33;
     memory[6832] = 32'd125;
     memory[6833] = 32'd156;
     memory[6834] = 32'd22;
     memory[6835] = 32'd102;
     memory[6836] = 32'd209;
     memory[6837] = 32'd98;
     memory[6838] = 32'd19;
     memory[6839] = 32'd0;
     memory[6840] = 32'd173;
     memory[6841] = 32'd173;
     memory[6842] = 32'd176;
     memory[6843] = 32'd81;
     memory[6844] = 32'd119;
     memory[6845] = 32'd22;
     memory[6846] = 32'd53;
     memory[6847] = 32'd182;
     memory[6848] = 32'd126;
     memory[6849] = 32'd88;
     memory[6850] = 32'd246;
     memory[6851] = 32'd148;
     memory[6852] = 32'd41;
     memory[6853] = 32'd133;
     memory[6854] = 32'd49;
     memory[6855] = 32'd94;
     memory[6856] = 32'd253;
     memory[6857] = 32'd180;
     memory[6858] = 32'd128;
     memory[6859] = 32'd212;
     memory[6860] = 32'd234;
     memory[6861] = 32'd144;
     memory[6862] = 32'd0;
     memory[6863] = 32'd211;
     memory[6864] = 32'd142;
     memory[6865] = 32'd68;
     memory[6866] = 32'd41;
     memory[6867] = 32'd79;
     memory[6868] = 32'd20;
     memory[6869] = 32'd90;
     memory[6870] = 32'd242;
     memory[6871] = 32'd218;
     memory[6872] = 32'd185;
     memory[6873] = 32'd219;
     memory[6874] = 32'd117;
     memory[6875] = 32'd78;
     memory[6876] = 32'd30;
     memory[6877] = 32'd29;
     memory[6878] = 32'd12;
     memory[6879] = 32'd120;
     memory[6880] = 32'd135;
     memory[6881] = 32'd188;
     memory[6882] = 32'd50;
     memory[6883] = 32'd125;
     memory[6884] = 32'd85;
     memory[6885] = 32'd143;
     memory[6886] = 32'd10;
     memory[6887] = 32'd22;
     memory[6888] = 32'd137;
     memory[6889] = 32'd158;
     memory[6890] = 32'd138;
     memory[6891] = 32'd50;
     memory[6892] = 32'd211;
     memory[6893] = 32'd229;
     memory[6894] = 32'd19;
     memory[6895] = 32'd40;
     memory[6896] = 32'd138;
     memory[6897] = 32'd119;
     memory[6898] = 32'd83;
     memory[6899] = 32'd212;
     memory[6900] = 32'd144;
     memory[6901] = 32'd4;
     memory[6902] = 32'd246;
     memory[6903] = 32'd153;
     memory[6904] = 32'd168;
     memory[6905] = 32'd254;
     memory[6906] = 32'd166;
     memory[6907] = 32'd57;
     memory[6908] = 32'd0;
     memory[6909] = 32'd188;
     memory[6910] = 32'd181;
     memory[6911] = 32'd248;
     memory[6912] = 32'd30;
     memory[6913] = 32'd217;
     memory[6914] = 32'd235;
     memory[6915] = 32'd26;
     memory[6916] = 32'd202;
     memory[6917] = 32'd11;
     memory[6918] = 32'd34;
     memory[6919] = 32'd110;
     memory[6920] = 32'd188;
     memory[6921] = 32'd204;
     memory[6922] = 32'd218;
     memory[6923] = 32'd253;
     memory[6924] = 32'd2;
     memory[6925] = 32'd99;
     memory[6926] = 32'd27;
     memory[6927] = 32'd202;
     memory[6928] = 32'd124;
     memory[6929] = 32'd25;
     memory[6930] = 32'd190;
     memory[6931] = 32'd75;
     memory[6932] = 32'd216;
     memory[6933] = 32'd144;
     memory[6934] = 32'd83;
     memory[6935] = 32'd216;
     memory[6936] = 32'd73;
     memory[6937] = 32'd152;
     memory[6938] = 32'd145;
     memory[6939] = 32'd2;
     memory[6940] = 32'd240;
     memory[6941] = 32'd2;
     memory[6942] = 32'd201;
     memory[6943] = 32'd16;
     memory[6944] = 32'd129;
     memory[6945] = 32'd173;
     memory[6946] = 32'd24;
     memory[6947] = 32'd11;
     memory[6948] = 32'd47;
     memory[6949] = 32'd73;
     memory[6950] = 32'd44;
     memory[6951] = 32'd36;
     memory[6952] = 32'd25;
     memory[6953] = 32'd239;
     memory[6954] = 32'd8;
     memory[6955] = 32'd151;
     memory[6956] = 32'd159;
     memory[6957] = 32'd159;
     memory[6958] = 32'd188;
     memory[6959] = 32'd191;
     memory[6960] = 32'd26;
     memory[6961] = 32'd11;
     memory[6962] = 32'd190;
     memory[6963] = 32'd182;
     memory[6964] = 32'd29;
     memory[6965] = 32'd161;
     memory[6966] = 32'd216;
     memory[6967] = 32'd196;
     memory[6968] = 32'd169;
     memory[6969] = 32'd21;
     memory[6970] = 32'd94;
     memory[6971] = 32'd248;
     memory[6972] = 32'd48;
     memory[6973] = 32'd209;
     memory[6974] = 32'd167;
     memory[6975] = 32'd199;
     memory[6976] = 32'd166;
     memory[6977] = 32'd186;
     memory[6978] = 32'd199;
     memory[6979] = 32'd235;
     memory[6980] = 32'd137;
     memory[6981] = 32'd49;
     memory[6982] = 32'd216;
     memory[6983] = 32'd199;
     memory[6984] = 32'd211;
     memory[6985] = 32'd93;
     memory[6986] = 32'd165;
     memory[6987] = 32'd95;
     memory[6988] = 32'd159;
     memory[6989] = 32'd150;
     memory[6990] = 32'd39;
     memory[6991] = 32'd27;
     memory[6992] = 32'd95;
     memory[6993] = 32'd244;
     memory[6994] = 32'd23;
     memory[6995] = 32'd54;
     memory[6996] = 32'd82;
     memory[6997] = 32'd18;
     memory[6998] = 32'd253;
     memory[6999] = 32'd24;
     memory[7000] = 32'd85;
     memory[7001] = 32'd25;
     memory[7002] = 32'd92;
     memory[7003] = 32'd183;
     memory[7004] = 32'd39;
     memory[7005] = 32'd113;
     memory[7006] = 32'd56;
     memory[7007] = 32'd251;
     memory[7008] = 32'd214;
     memory[7009] = 32'd180;
     memory[7010] = 32'd124;
     memory[7011] = 32'd251;
     memory[7012] = 32'd145;
     memory[7013] = 32'd101;
     memory[7014] = 32'd150;
     memory[7015] = 32'd160;
     memory[7016] = 32'd212;
     memory[7017] = 32'd11;
     memory[7018] = 32'd56;
     memory[7019] = 32'd175;
     memory[7020] = 32'd208;
     memory[7021] = 32'd126;
     memory[7022] = 32'd202;
     memory[7023] = 32'd153;
     memory[7024] = 32'd228;
     memory[7025] = 32'd170;
     memory[7026] = 32'd86;
     memory[7027] = 32'd192;
     memory[7028] = 32'd185;
     memory[7029] = 32'd22;
     memory[7030] = 32'd86;
     memory[7031] = 32'd205;
     memory[7032] = 32'd102;
     memory[7033] = 32'd104;
     memory[7034] = 32'd208;
     memory[7035] = 32'd166;
     memory[7036] = 32'd26;
     memory[7037] = 32'd118;
     memory[7038] = 32'd208;
     memory[7039] = 32'd99;
     memory[7040] = 32'd64;
     memory[7041] = 32'd41;
     memory[7042] = 32'd16;
     memory[7043] = 32'd77;
     memory[7044] = 32'd230;
     memory[7045] = 32'd61;
     memory[7046] = 32'd195;
     memory[7047] = 32'd35;
     memory[7048] = 32'd66;
     memory[7049] = 32'd151;
     memory[7050] = 32'd7;
     memory[7051] = 32'd80;
     memory[7052] = 32'd51;
     memory[7053] = 32'd140;
     memory[7054] = 32'd18;
     memory[7055] = 32'd86;
     memory[7056] = 32'd181;
     memory[7057] = 32'd217;
     memory[7058] = 32'd115;
     memory[7059] = 32'd220;
     memory[7060] = 32'd194;
     memory[7061] = 32'd129;
     memory[7062] = 32'd245;
     memory[7063] = 32'd13;
     memory[7064] = 32'd115;
     memory[7065] = 32'd219;
     memory[7066] = 32'd128;
     memory[7067] = 32'd208;
     memory[7068] = 32'd39;
     memory[7069] = 32'd175;
     memory[7070] = 32'd72;
     memory[7071] = 32'd182;
     memory[7072] = 32'd101;
     memory[7073] = 32'd41;
     memory[7074] = 32'd196;
     memory[7075] = 32'd198;
     memory[7076] = 32'd245;
     memory[7077] = 32'd86;
     memory[7078] = 32'd252;
     memory[7079] = 32'd88;
     memory[7080] = 32'd164;
     memory[7081] = 32'd152;
     memory[7082] = 32'd119;
     memory[7083] = 32'd133;
     memory[7084] = 32'd145;
     memory[7085] = 32'd149;
     memory[7086] = 32'd34;
     memory[7087] = 32'd40;
     memory[7088] = 32'd113;
     memory[7089] = 32'd178;
     memory[7090] = 32'd32;
     memory[7091] = 32'd129;
     memory[7092] = 32'd17;
     memory[7093] = 32'd184;
     memory[7094] = 32'd90;
     memory[7095] = 32'd28;
     memory[7096] = 32'd6;
     memory[7097] = 32'd97;
     memory[7098] = 32'd7;
     memory[7099] = 32'd126;
     memory[7100] = 32'd129;
     memory[7101] = 32'd251;
     memory[7102] = 32'd5;
     memory[7103] = 32'd194;
     memory[7104] = 32'd57;
     memory[7105] = 32'd59;
     memory[7106] = 32'd127;
     memory[7107] = 32'd82;
     memory[7108] = 32'd159;
     memory[7109] = 32'd74;
     memory[7110] = 32'd193;
     memory[7111] = 32'd151;
     memory[7112] = 32'd202;
     memory[7113] = 32'd172;
     memory[7114] = 32'd152;
     memory[7115] = 32'd243;
     memory[7116] = 32'd247;
     memory[7117] = 32'd182;
     memory[7118] = 32'd245;
     memory[7119] = 32'd84;
     memory[7120] = 32'd199;
     memory[7121] = 32'd215;
     memory[7122] = 32'd122;
     memory[7123] = 32'd95;
     memory[7124] = 32'd8;
     memory[7125] = 32'd98;
     memory[7126] = 32'd235;
     memory[7127] = 32'd177;
     memory[7128] = 32'd57;
     memory[7129] = 32'd124;
     memory[7130] = 32'd32;
     memory[7131] = 32'd247;
     memory[7132] = 32'd200;
     memory[7133] = 32'd134;
     memory[7134] = 32'd58;
     memory[7135] = 32'd130;
     memory[7136] = 32'd141;
     memory[7137] = 32'd76;
     memory[7138] = 32'd25;
     memory[7139] = 32'd226;
     memory[7140] = 32'd174;
     memory[7141] = 32'd188;
     memory[7142] = 32'd233;
     memory[7143] = 32'd80;
     memory[7144] = 32'd170;
     memory[7145] = 32'd181;
     memory[7146] = 32'd119;
     memory[7147] = 32'd116;
     memory[7148] = 32'd140;
     memory[7149] = 32'd184;
     memory[7150] = 32'd217;
     memory[7151] = 32'd198;
     memory[7152] = 32'd17;
     memory[7153] = 32'd105;
     memory[7154] = 32'd76;
     memory[7155] = 32'd130;
     memory[7156] = 32'd218;
     memory[7157] = 32'd109;
     memory[7158] = 32'd145;
     memory[7159] = 32'd92;
     memory[7160] = 32'd144;
     memory[7161] = 32'd172;
     memory[7162] = 32'd107;
     memory[7163] = 32'd173;
     memory[7164] = 32'd79;
     memory[7165] = 32'd105;
     memory[7166] = 32'd28;
     memory[7167] = 32'd46;
     memory[7168] = 32'd209;
     memory[7169] = 32'd182;
     memory[7170] = 32'd182;
     memory[7171] = 32'd225;
     memory[7172] = 32'd215;
     memory[7173] = 32'd17;
     memory[7174] = 32'd79;
     memory[7175] = 32'd224;
     memory[7176] = 32'd180;
     memory[7177] = 32'd191;
     memory[7178] = 32'd198;
     memory[7179] = 32'd5;
     memory[7180] = 32'd222;
     memory[7181] = 32'd197;
     memory[7182] = 32'd36;
     memory[7183] = 32'd43;
     memory[7184] = 32'd14;
     memory[7185] = 32'd131;
     memory[7186] = 32'd242;
     memory[7187] = 32'd3;
     memory[7188] = 32'd118;
     memory[7189] = 32'd218;
     memory[7190] = 32'd226;
     memory[7191] = 32'd206;
     memory[7192] = 32'd14;
     memory[7193] = 32'd235;
     memory[7194] = 32'd27;
     memory[7195] = 32'd139;
     memory[7196] = 32'd99;
     memory[7197] = 32'd148;
     memory[7198] = 32'd188;
     memory[7199] = 32'd13;
     memory[7200] = 32'd24;
     memory[7201] = 32'd180;
     memory[7202] = 32'd160;
     memory[7203] = 32'd223;
     memory[7204] = 32'd149;
     memory[7205] = 32'd65;
     memory[7206] = 32'd54;
     memory[7207] = 32'd242;
     memory[7208] = 32'd226;
     memory[7209] = 32'd38;
     memory[7210] = 32'd168;
     memory[7211] = 32'd76;
     memory[7212] = 32'd176;
     memory[7213] = 32'd136;
     memory[7214] = 32'd154;
     memory[7215] = 32'd206;
     memory[7216] = 32'd2;
     memory[7217] = 32'd15;
     memory[7218] = 32'd74;
     memory[7219] = 32'd180;
     memory[7220] = 32'd49;
     memory[7221] = 32'd207;
     memory[7222] = 32'd22;
     memory[7223] = 32'd253;
     memory[7224] = 32'd141;
     memory[7225] = 32'd200;
     memory[7226] = 32'd151;
     memory[7227] = 32'd149;
     memory[7228] = 32'd14;
     memory[7229] = 32'd205;
     memory[7230] = 32'd54;
     memory[7231] = 32'd143;
     memory[7232] = 32'd220;
     memory[7233] = 32'd157;
     memory[7234] = 32'd126;
     memory[7235] = 32'd45;
     memory[7236] = 32'd244;
     memory[7237] = 32'd103;
     memory[7238] = 32'd21;
     memory[7239] = 32'd194;
     memory[7240] = 32'd33;
     memory[7241] = 32'd42;
     memory[7242] = 32'd181;
     memory[7243] = 32'd1;
     memory[7244] = 32'd127;
     memory[7245] = 32'd68;
     memory[7246] = 32'd110;
     memory[7247] = 32'd181;
     memory[7248] = 32'd132;
     memory[7249] = 32'd184;
     memory[7250] = 32'd160;
     memory[7251] = 32'd48;
     memory[7252] = 32'd227;
     memory[7253] = 32'd30;
     memory[7254] = 32'd205;
     memory[7255] = 32'd140;
     memory[7256] = 32'd218;
     memory[7257] = 32'd9;
     memory[7258] = 32'd37;
     memory[7259] = 32'd6;
     memory[7260] = 32'd209;
     memory[7261] = 32'd127;
     memory[7262] = 32'd43;
     memory[7263] = 32'd158;
     memory[7264] = 32'd132;
     memory[7265] = 32'd213;
     memory[7266] = 32'd123;
     memory[7267] = 32'd248;
     memory[7268] = 32'd134;
     memory[7269] = 32'd7;
     memory[7270] = 32'd71;
     memory[7271] = 32'd198;
     memory[7272] = 32'd140;
     memory[7273] = 32'd140;
     memory[7274] = 32'd93;
     memory[7275] = 32'd72;
     memory[7276] = 32'd143;
     memory[7277] = 32'd0;
     memory[7278] = 32'd223;
     memory[7279] = 32'd165;
     memory[7280] = 32'd155;
     memory[7281] = 32'd95;
     memory[7282] = 32'd191;
     memory[7283] = 32'd145;
     memory[7284] = 32'd161;
     memory[7285] = 32'd161;
     memory[7286] = 32'd243;
     memory[7287] = 32'd210;
     memory[7288] = 32'd223;
     memory[7289] = 32'd236;
     memory[7290] = 32'd245;
     memory[7291] = 32'd102;
     memory[7292] = 32'd185;
     memory[7293] = 32'd14;
     memory[7294] = 32'd45;
     memory[7295] = 32'd129;
     memory[7296] = 32'd244;
     memory[7297] = 32'd107;
     memory[7298] = 32'd206;
     memory[7299] = 32'd249;
     memory[7300] = 32'd180;
     memory[7301] = 32'd5;
     memory[7302] = 32'd50;
     memory[7303] = 32'd208;
     memory[7304] = 32'd119;
     memory[7305] = 32'd93;
     memory[7306] = 32'd145;
     memory[7307] = 32'd218;
     memory[7308] = 32'd233;
     memory[7309] = 32'd11;
     memory[7310] = 32'd29;
     memory[7311] = 32'd24;
     memory[7312] = 32'd206;
     memory[7313] = 32'd53;
     memory[7314] = 32'd132;
     memory[7315] = 32'd81;
     memory[7316] = 32'd45;
     memory[7317] = 32'd219;
     memory[7318] = 32'd251;
     memory[7319] = 32'd252;
     memory[7320] = 32'd115;
     memory[7321] = 32'd113;
     memory[7322] = 32'd48;
     memory[7323] = 32'd141;
     memory[7324] = 32'd53;
     memory[7325] = 32'd78;
     memory[7326] = 32'd232;
     memory[7327] = 32'd126;
     memory[7328] = 32'd206;
     memory[7329] = 32'd237;
     memory[7330] = 32'd171;
     memory[7331] = 32'd139;
     memory[7332] = 32'd142;
     memory[7333] = 32'd75;
     memory[7334] = 32'd70;
     memory[7335] = 32'd76;
     memory[7336] = 32'd73;
     memory[7337] = 32'd42;
     memory[7338] = 32'd154;
     memory[7339] = 32'd245;
     memory[7340] = 32'd185;
     memory[7341] = 32'd248;
     memory[7342] = 32'd38;
     memory[7343] = 32'd194;
     memory[7344] = 32'd89;
     memory[7345] = 32'd9;
     memory[7346] = 32'd72;
     memory[7347] = 32'd190;
     memory[7348] = 32'd108;
     memory[7349] = 32'd125;
     memory[7350] = 32'd247;
     memory[7351] = 32'd211;
     memory[7352] = 32'd246;
     memory[7353] = 32'd171;
     memory[7354] = 32'd185;
     memory[7355] = 32'd253;
     memory[7356] = 32'd71;
     memory[7357] = 32'd115;
     memory[7358] = 32'd37;
     memory[7359] = 32'd7;
     memory[7360] = 32'd10;
     memory[7361] = 32'd143;
     memory[7362] = 32'd131;
     memory[7363] = 32'd94;
     memory[7364] = 32'd186;
     memory[7365] = 32'd75;
     memory[7366] = 32'd18;
     memory[7367] = 32'd72;
     memory[7368] = 32'd191;
     memory[7369] = 32'd244;
     memory[7370] = 32'd9;
     memory[7371] = 32'd119;
     memory[7372] = 32'd39;
     memory[7373] = 32'd163;
     memory[7374] = 32'd165;
     memory[7375] = 32'd119;
     memory[7376] = 32'd144;
     memory[7377] = 32'd198;
     memory[7378] = 32'd79;
     memory[7379] = 32'd227;
     memory[7380] = 32'd116;
     memory[7381] = 32'd60;
     memory[7382] = 32'd134;
     memory[7383] = 32'd55;
     memory[7384] = 32'd171;
     memory[7385] = 32'd134;
     memory[7386] = 32'd192;
     memory[7387] = 32'd249;
     memory[7388] = 32'd247;
     memory[7389] = 32'd60;
     memory[7390] = 32'd104;
     memory[7391] = 32'd250;
     memory[7392] = 32'd158;
     memory[7393] = 32'd237;
     memory[7394] = 32'd41;
     memory[7395] = 32'd247;
     memory[7396] = 32'd158;
     memory[7397] = 32'd19;
     memory[7398] = 32'd161;
     memory[7399] = 32'd143;
     memory[7400] = 32'd93;
     memory[7401] = 32'd191;
     memory[7402] = 32'd60;
     memory[7403] = 32'd171;
     memory[7404] = 32'd179;
     memory[7405] = 32'd60;
     memory[7406] = 32'd19;
     memory[7407] = 32'd47;
     memory[7408] = 32'd164;
     memory[7409] = 32'd128;
     memory[7410] = 32'd196;
     memory[7411] = 32'd201;
     memory[7412] = 32'd188;
     memory[7413] = 32'd201;
     memory[7414] = 32'd105;
     memory[7415] = 32'd28;
     memory[7416] = 32'd136;
     memory[7417] = 32'd253;
     memory[7418] = 32'd58;
     memory[7419] = 32'd181;
     memory[7420] = 32'd216;
     memory[7421] = 32'd60;
     memory[7422] = 32'd147;
     memory[7423] = 32'd78;
     memory[7424] = 32'd35;
     memory[7425] = 32'd107;
     memory[7426] = 32'd188;
     memory[7427] = 32'd223;
     memory[7428] = 32'd240;
     memory[7429] = 32'd142;
     memory[7430] = 32'd26;
     memory[7431] = 32'd193;
     memory[7432] = 32'd242;
     memory[7433] = 32'd55;
     memory[7434] = 32'd2;
     memory[7435] = 32'd184;
     memory[7436] = 32'd182;
     memory[7437] = 32'd222;
     memory[7438] = 32'd250;
     memory[7439] = 32'd96;
     memory[7440] = 32'd215;
     memory[7441] = 32'd132;
     memory[7442] = 32'd193;
     memory[7443] = 32'd110;
     memory[7444] = 32'd30;
     memory[7445] = 32'd56;
     memory[7446] = 32'd146;
     memory[7447] = 32'd68;
     memory[7448] = 32'd129;
     memory[7449] = 32'd85;
     memory[7450] = 32'd183;
     memory[7451] = 32'd64;
     memory[7452] = 32'd185;
     memory[7453] = 32'd5;
     memory[7454] = 32'd55;
     memory[7455] = 32'd191;
     memory[7456] = 32'd120;
     memory[7457] = 32'd190;
     memory[7458] = 32'd121;
     memory[7459] = 32'd128;
     memory[7460] = 32'd137;
     memory[7461] = 32'd127;
     memory[7462] = 32'd214;
     memory[7463] = 32'd6;
     memory[7464] = 32'd53;
     memory[7465] = 32'd243;
     memory[7466] = 32'd235;
     memory[7467] = 32'd25;
     memory[7468] = 32'd11;
     memory[7469] = 32'd95;
     memory[7470] = 32'd193;
     memory[7471] = 32'd12;
     memory[7472] = 32'd49;
     memory[7473] = 32'd121;
     memory[7474] = 32'd222;
     memory[7475] = 32'd16;
     memory[7476] = 32'd10;
     memory[7477] = 32'd5;
     memory[7478] = 32'd95;
     memory[7479] = 32'd219;
     memory[7480] = 32'd173;
     memory[7481] = 32'd146;
     memory[7482] = 32'd74;
     memory[7483] = 32'd81;
     memory[7484] = 32'd3;
     memory[7485] = 32'd36;
     memory[7486] = 32'd101;
     memory[7487] = 32'd65;
     memory[7488] = 32'd220;
     memory[7489] = 32'd2;
     memory[7490] = 32'd49;
     memory[7491] = 32'd230;
     memory[7492] = 32'd30;
     memory[7493] = 32'd78;
     memory[7494] = 32'd138;
     memory[7495] = 32'd119;
     memory[7496] = 32'd108;
     memory[7497] = 32'd55;
     memory[7498] = 32'd157;
     memory[7499] = 32'd196;
     memory[7500] = 32'd101;
     memory[7501] = 32'd202;
     memory[7502] = 32'd99;
     memory[7503] = 32'd195;
     memory[7504] = 32'd248;
     memory[7505] = 32'd94;
     memory[7506] = 32'd71;
     memory[7507] = 32'd1;
     memory[7508] = 32'd132;
     memory[7509] = 32'd250;
     memory[7510] = 32'd148;
     memory[7511] = 32'd85;
     memory[7512] = 32'd114;
     memory[7513] = 32'd215;
     memory[7514] = 32'd124;
     memory[7515] = 32'd136;
     memory[7516] = 32'd136;
     memory[7517] = 32'd8;
     memory[7518] = 32'd156;
     memory[7519] = 32'd81;
     memory[7520] = 32'd186;
     memory[7521] = 32'd219;
     memory[7522] = 32'd117;
     memory[7523] = 32'd196;
     memory[7524] = 32'd183;
     memory[7525] = 32'd38;
     memory[7526] = 32'd169;
     memory[7527] = 32'd12;
     memory[7528] = 32'd55;
     memory[7529] = 32'd115;
     memory[7530] = 32'd159;
     memory[7531] = 32'd49;
     memory[7532] = 32'd156;
     memory[7533] = 32'd142;
     memory[7534] = 32'd106;
     memory[7535] = 32'd80;
     memory[7536] = 32'd117;
     memory[7537] = 32'd5;
     memory[7538] = 32'd28;
     memory[7539] = 32'd11;
     memory[7540] = 32'd196;
     memory[7541] = 32'd175;
     memory[7542] = 32'd53;
     memory[7543] = 32'd138;
     memory[7544] = 32'd211;
     memory[7545] = 32'd95;
     memory[7546] = 32'd164;
     memory[7547] = 32'd4;
     memory[7548] = 32'd250;
     memory[7549] = 32'd79;
     memory[7550] = 32'd183;
     memory[7551] = 32'd187;
     memory[7552] = 32'd11;
     memory[7553] = 32'd132;
     memory[7554] = 32'd133;
     memory[7555] = 32'd206;
     memory[7556] = 32'd186;
     memory[7557] = 32'd220;
     memory[7558] = 32'd120;
     memory[7559] = 32'd21;
     memory[7560] = 32'd50;
     memory[7561] = 32'd244;
     memory[7562] = 32'd177;
     memory[7563] = 32'd183;
     memory[7564] = 32'd241;
     memory[7565] = 32'd233;
     memory[7566] = 32'd20;
     memory[7567] = 32'd31;
     memory[7568] = 32'd185;
     memory[7569] = 32'd201;
     memory[7570] = 32'd25;
     memory[7571] = 32'd74;
     memory[7572] = 32'd103;
     memory[7573] = 32'd157;
     memory[7574] = 32'd217;
     memory[7575] = 32'd189;
     memory[7576] = 32'd245;
     memory[7577] = 32'd204;
     memory[7578] = 32'd46;
     memory[7579] = 32'd166;
     memory[7580] = 32'd126;
     memory[7581] = 32'd91;
     memory[7582] = 32'd32;
     memory[7583] = 32'd202;
     memory[7584] = 32'd31;
     memory[7585] = 32'd197;
     memory[7586] = 32'd92;
     memory[7587] = 32'd168;
     memory[7588] = 32'd156;
     memory[7589] = 32'd185;
     memory[7590] = 32'd91;
     memory[7591] = 32'd63;
     memory[7592] = 32'd126;
     memory[7593] = 32'd181;
     memory[7594] = 32'd78;
     memory[7595] = 32'd49;
     memory[7596] = 32'd201;
     memory[7597] = 32'd212;
     memory[7598] = 32'd50;
     memory[7599] = 32'd28;
     memory[7600] = 32'd151;
     memory[7601] = 32'd106;
     memory[7602] = 32'd0;
     memory[7603] = 32'd104;
     memory[7604] = 32'd24;
     memory[7605] = 32'd35;
     memory[7606] = 32'd89;
     memory[7607] = 32'd227;
     memory[7608] = 32'd227;
     memory[7609] = 32'd238;
     memory[7610] = 32'd151;
     memory[7611] = 32'd107;
     memory[7612] = 32'd56;
     memory[7613] = 32'd14;
     memory[7614] = 32'd49;
     memory[7615] = 32'd229;
     memory[7616] = 32'd121;
     memory[7617] = 32'd154;
     memory[7618] = 32'd41;
     memory[7619] = 32'd3;
     memory[7620] = 32'd155;
     memory[7621] = 32'd0;
     memory[7622] = 32'd123;
     memory[7623] = 32'd20;
     memory[7624] = 32'd50;
     memory[7625] = 32'd25;
     memory[7626] = 32'd4;
     memory[7627] = 32'd164;
     memory[7628] = 32'd134;
     memory[7629] = 32'd171;
     memory[7630] = 32'd150;
     memory[7631] = 32'd72;
     memory[7632] = 32'd117;
     memory[7633] = 32'd183;
     memory[7634] = 32'd226;
     memory[7635] = 32'd191;
     memory[7636] = 32'd104;
     memory[7637] = 32'd217;
     memory[7638] = 32'd165;
     memory[7639] = 32'd238;
     memory[7640] = 32'd67;
     memory[7641] = 32'd202;
     memory[7642] = 32'd168;
     memory[7643] = 32'd110;
     memory[7644] = 32'd197;
     memory[7645] = 32'd16;
     memory[7646] = 32'd167;
     memory[7647] = 32'd25;
     memory[7648] = 32'd227;
     memory[7649] = 32'd190;
     memory[7650] = 32'd218;
     memory[7651] = 32'd64;
     memory[7652] = 32'd158;
     memory[7653] = 32'd66;
     memory[7654] = 32'd3;
     memory[7655] = 32'd129;
     memory[7656] = 32'd169;
     memory[7657] = 32'd49;
     memory[7658] = 32'd71;
     memory[7659] = 32'd34;
     memory[7660] = 32'd218;
     memory[7661] = 32'd137;
     memory[7662] = 32'd244;
     memory[7663] = 32'd16;
     memory[7664] = 32'd42;
     memory[7665] = 32'd124;
     memory[7666] = 32'd71;
     memory[7667] = 32'd221;
     memory[7668] = 32'd150;
     memory[7669] = 32'd48;
     memory[7670] = 32'd7;
     memory[7671] = 32'd239;
     memory[7672] = 32'd183;
     memory[7673] = 32'd165;
     memory[7674] = 32'd26;
     memory[7675] = 32'd73;
     memory[7676] = 32'd251;
     memory[7677] = 32'd26;
     memory[7678] = 32'd67;
     memory[7679] = 32'd64;
     memory[7680] = 32'd50;
     memory[7681] = 32'd96;
     memory[7682] = 32'd61;
     memory[7683] = 32'd136;
     memory[7684] = 32'd220;
     memory[7685] = 32'd183;
     memory[7686] = 32'd252;
     memory[7687] = 32'd59;
     memory[7688] = 32'd222;
     memory[7689] = 32'd189;
     memory[7690] = 32'd135;
     memory[7691] = 32'd76;
     memory[7692] = 32'd34;
     memory[7693] = 32'd245;
     memory[7694] = 32'd230;
     memory[7695] = 32'd223;
     memory[7696] = 32'd240;
     memory[7697] = 32'd58;
     memory[7698] = 32'd73;
     memory[7699] = 32'd231;
     memory[7700] = 32'd105;
     memory[7701] = 32'd48;
     memory[7702] = 32'd114;
     memory[7703] = 32'd167;
     memory[7704] = 32'd155;
     memory[7705] = 32'd201;
     memory[7706] = 32'd235;
     memory[7707] = 32'd25;
     memory[7708] = 32'd190;
     memory[7709] = 32'd177;
     memory[7710] = 32'd252;
     memory[7711] = 32'd64;
     memory[7712] = 32'd106;
     memory[7713] = 32'd242;
     memory[7714] = 32'd210;
     memory[7715] = 32'd86;
     memory[7716] = 32'd164;
     memory[7717] = 32'd25;
     memory[7718] = 32'd112;
     memory[7719] = 32'd40;
     memory[7720] = 32'd163;
     memory[7721] = 32'd24;
     memory[7722] = 32'd242;
     memory[7723] = 32'd223;
     memory[7724] = 32'd212;
     memory[7725] = 32'd157;
     memory[7726] = 32'd222;
     memory[7727] = 32'd164;
     memory[7728] = 32'd59;
     memory[7729] = 32'd37;
     memory[7730] = 32'd20;
     memory[7731] = 32'd127;
     memory[7732] = 32'd173;
     memory[7733] = 32'd78;
     memory[7734] = 32'd203;
     memory[7735] = 32'd181;
     memory[7736] = 32'd105;
     memory[7737] = 32'd80;
     memory[7738] = 32'd97;
     memory[7739] = 32'd203;
     memory[7740] = 32'd215;
     memory[7741] = 32'd181;
     memory[7742] = 32'd198;
     memory[7743] = 32'd149;
     memory[7744] = 32'd12;
     memory[7745] = 32'd138;
     memory[7746] = 32'd123;
     memory[7747] = 32'd5;
     memory[7748] = 32'd0;
     memory[7749] = 32'd188;
     memory[7750] = 32'd21;
     memory[7751] = 32'd126;
     memory[7752] = 32'd11;
     memory[7753] = 32'd36;
     memory[7754] = 32'd107;
     memory[7755] = 32'd51;
     memory[7756] = 32'd34;
     memory[7757] = 32'd254;
     memory[7758] = 32'd59;
     memory[7759] = 32'd165;
     memory[7760] = 32'd81;
     memory[7761] = 32'd57;
     memory[7762] = 32'd29;
     memory[7763] = 32'd73;
     memory[7764] = 32'd62;
     memory[7765] = 32'd63;
     memory[7766] = 32'd74;
     memory[7767] = 32'd190;
     memory[7768] = 32'd75;
     memory[7769] = 32'd134;
     memory[7770] = 32'd254;
     memory[7771] = 32'd67;
     memory[7772] = 32'd157;
     memory[7773] = 32'd145;
     memory[7774] = 32'd228;
     memory[7775] = 32'd192;
     memory[7776] = 32'd99;
     memory[7777] = 32'd93;
     memory[7778] = 32'd158;
     memory[7779] = 32'd24;
     memory[7780] = 32'd247;
     memory[7781] = 32'd238;
     memory[7782] = 32'd222;
     memory[7783] = 32'd17;
     memory[7784] = 32'd84;
     memory[7785] = 32'd71;
     memory[7786] = 32'd139;
     memory[7787] = 32'd28;
     memory[7788] = 32'd35;
     memory[7789] = 32'd18;
     memory[7790] = 32'd71;
     memory[7791] = 32'd118;
     memory[7792] = 32'd168;
     memory[7793] = 32'd212;
     memory[7794] = 32'd230;
     memory[7795] = 32'd124;
     memory[7796] = 32'd14;
     memory[7797] = 32'd82;
     memory[7798] = 32'd166;
     memory[7799] = 32'd137;
     memory[7800] = 32'd241;
     memory[7801] = 32'd68;
     memory[7802] = 32'd145;
     memory[7803] = 32'd192;
     memory[7804] = 32'd107;
     memory[7805] = 32'd101;
     memory[7806] = 32'd135;
     memory[7807] = 32'd117;
     memory[7808] = 32'd66;
     memory[7809] = 32'd200;
     memory[7810] = 32'd171;
     memory[7811] = 32'd167;
     memory[7812] = 32'd155;
     memory[7813] = 32'd21;
     memory[7814] = 32'd24;
     memory[7815] = 32'd136;
     memory[7816] = 32'd169;
     memory[7817] = 32'd203;
     memory[7818] = 32'd137;
     memory[7819] = 32'd123;
     memory[7820] = 32'd174;
     memory[7821] = 32'd253;
     memory[7822] = 32'd80;
     memory[7823] = 32'd211;
     memory[7824] = 32'd174;
     memory[7825] = 32'd186;
     memory[7826] = 32'd116;
     memory[7827] = 32'd111;
     memory[7828] = 32'd125;
     memory[7829] = 32'd73;
     memory[7830] = 32'd19;
     memory[7831] = 32'd235;
     memory[7832] = 32'd245;
     memory[7833] = 32'd42;
     memory[7834] = 32'd129;
     memory[7835] = 32'd36;
     memory[7836] = 32'd228;
     memory[7837] = 32'd65;
     memory[7838] = 32'd194;
     memory[7839] = 32'd210;
     memory[7840] = 32'd137;
     memory[7841] = 32'd242;
     memory[7842] = 32'd122;
     memory[7843] = 32'd178;
     memory[7844] = 32'd171;
     memory[7845] = 32'd191;
     memory[7846] = 32'd22;
     memory[7847] = 32'd252;
     memory[7848] = 32'd149;
     memory[7849] = 32'd52;
     memory[7850] = 32'd253;
     memory[7851] = 32'd153;
     memory[7852] = 32'd212;
     memory[7853] = 32'd244;
     memory[7854] = 32'd196;
     memory[7855] = 32'd48;
     memory[7856] = 32'd226;
     memory[7857] = 32'd29;
     memory[7858] = 32'd108;
     memory[7859] = 32'd88;
     memory[7860] = 32'd1;
     memory[7861] = 32'd15;
     memory[7862] = 32'd97;
     memory[7863] = 32'd187;
     memory[7864] = 32'd176;
     memory[7865] = 32'd12;
     memory[7866] = 32'd81;
     memory[7867] = 32'd114;
     memory[7868] = 32'd61;
     memory[7869] = 32'd150;
     memory[7870] = 32'd217;
     memory[7871] = 32'd151;
     memory[7872] = 32'd66;
     memory[7873] = 32'd168;
     memory[7874] = 32'd29;
     memory[7875] = 32'd149;
     memory[7876] = 32'd112;
     memory[7877] = 32'd151;
     memory[7878] = 32'd246;
     memory[7879] = 32'd72;
     memory[7880] = 32'd77;
     memory[7881] = 32'd246;
     memory[7882] = 32'd121;
     memory[7883] = 32'd44;
     memory[7884] = 32'd197;
     memory[7885] = 32'd183;
     memory[7886] = 32'd173;
     memory[7887] = 32'd19;
     memory[7888] = 32'd101;
     memory[7889] = 32'd79;
     memory[7890] = 32'd111;
     memory[7891] = 32'd182;
     memory[7892] = 32'd234;
     memory[7893] = 32'd165;
     memory[7894] = 32'd169;
     memory[7895] = 32'd197;
     memory[7896] = 32'd82;
     memory[7897] = 32'd121;
     memory[7898] = 32'd237;
     memory[7899] = 32'd236;
     memory[7900] = 32'd73;
     memory[7901] = 32'd14;
     memory[7902] = 32'd106;
     memory[7903] = 32'd243;
     memory[7904] = 32'd163;
     memory[7905] = 32'd38;
     memory[7906] = 32'd118;
     memory[7907] = 32'd219;
     memory[7908] = 32'd90;
     memory[7909] = 32'd206;
     memory[7910] = 32'd12;
     memory[7911] = 32'd110;
     memory[7912] = 32'd92;
     memory[7913] = 32'd187;
     memory[7914] = 32'd168;
     memory[7915] = 32'd172;
     memory[7916] = 32'd112;
     memory[7917] = 32'd182;
     memory[7918] = 32'd61;
     memory[7919] = 32'd130;
     memory[7920] = 32'd2;
     memory[7921] = 32'd192;
     memory[7922] = 32'd121;
     memory[7923] = 32'd47;
     memory[7924] = 32'd224;
     memory[7925] = 32'd142;
     memory[7926] = 32'd68;
     memory[7927] = 32'd14;
     memory[7928] = 32'd148;
     memory[7929] = 32'd73;
     memory[7930] = 32'd45;
     memory[7931] = 32'd189;
     memory[7932] = 32'd231;
     memory[7933] = 32'd167;
     memory[7934] = 32'd231;
     memory[7935] = 32'd143;
     memory[7936] = 32'd66;
     memory[7937] = 32'd44;
     memory[7938] = 32'd53;
     memory[7939] = 32'd24;
     memory[7940] = 32'd224;
     memory[7941] = 32'd52;
     memory[7942] = 32'd17;
     memory[7943] = 32'd86;
     memory[7944] = 32'd46;
     memory[7945] = 32'd128;
     memory[7946] = 32'd43;
     memory[7947] = 32'd163;
     memory[7948] = 32'd221;
     memory[7949] = 32'd66;
     memory[7950] = 32'd52;
     memory[7951] = 32'd167;
     memory[7952] = 32'd123;
     memory[7953] = 32'd83;
     memory[7954] = 32'd120;
     memory[7955] = 32'd49;
     memory[7956] = 32'd79;
     memory[7957] = 32'd159;
     memory[7958] = 32'd47;
     memory[7959] = 32'd4;
     memory[7960] = 32'd173;
     memory[7961] = 32'd41;
     memory[7962] = 32'd208;
     memory[7963] = 32'd230;
     memory[7964] = 32'd218;
     memory[7965] = 32'd129;
     memory[7966] = 32'd80;
     memory[7967] = 32'd24;
     memory[7968] = 32'd102;
     memory[7969] = 32'd95;
     memory[7970] = 32'd5;
     memory[7971] = 32'd190;
     memory[7972] = 32'd90;
     memory[7973] = 32'd27;
     memory[7974] = 32'd176;
     memory[7975] = 32'd199;
     memory[7976] = 32'd98;
     memory[7977] = 32'd173;
     memory[7978] = 32'd29;
     memory[7979] = 32'd96;
     memory[7980] = 32'd12;
     memory[7981] = 32'd99;
     memory[7982] = 32'd56;
     memory[7983] = 32'd206;
     memory[7984] = 32'd235;
     memory[7985] = 32'd174;
     memory[7986] = 32'd22;
     memory[7987] = 32'd124;
     memory[7988] = 32'd160;
     memory[7989] = 32'd100;
     memory[7990] = 32'd196;
     memory[7991] = 32'd124;
     memory[7992] = 32'd118;
     memory[7993] = 32'd195;
     memory[7994] = 32'd252;
     memory[7995] = 32'd11;
     memory[7996] = 32'd215;
     memory[7997] = 32'd53;
     memory[7998] = 32'd122;
     memory[7999] = 32'd18;
     memory[8000] = 32'd206;
     memory[8001] = 32'd42;
     memory[8002] = 32'd68;
     memory[8003] = 32'd194;
     memory[8004] = 32'd134;
     memory[8005] = 32'd137;
     memory[8006] = 32'd193;
     memory[8007] = 32'd86;
     memory[8008] = 32'd207;
     memory[8009] = 32'd111;
     memory[8010] = 32'd27;
     memory[8011] = 32'd15;
     memory[8012] = 32'd164;
     memory[8013] = 32'd29;
     memory[8014] = 32'd181;
     memory[8015] = 32'd235;
     memory[8016] = 32'd9;
     memory[8017] = 32'd142;
     memory[8018] = 32'd96;
     memory[8019] = 32'd181;
     memory[8020] = 32'd142;
     memory[8021] = 32'd180;
     memory[8022] = 32'd54;
     memory[8023] = 32'd74;
     memory[8024] = 32'd140;
     memory[8025] = 32'd90;
     memory[8026] = 32'd214;
     memory[8027] = 32'd216;
     memory[8028] = 32'd64;
     memory[8029] = 32'd105;
     memory[8030] = 32'd176;
     memory[8031] = 32'd243;
     memory[8032] = 32'd99;
     memory[8033] = 32'd197;
     memory[8034] = 32'd85;
     memory[8035] = 32'd100;
     memory[8036] = 32'd230;
     memory[8037] = 32'd22;
     memory[8038] = 32'd170;
     memory[8039] = 32'd140;
     memory[8040] = 32'd139;
     memory[8041] = 32'd58;
     memory[8042] = 32'd80;
     memory[8043] = 32'd157;
     memory[8044] = 32'd146;
     memory[8045] = 32'd136;
     memory[8046] = 32'd6;
     memory[8047] = 32'd241;
     memory[8048] = 32'd10;
     memory[8049] = 32'd106;
     memory[8050] = 32'd114;
     memory[8051] = 32'd84;
     memory[8052] = 32'd244;
     memory[8053] = 32'd140;
     memory[8054] = 32'd68;
     memory[8055] = 32'd139;
     memory[8056] = 32'd135;
     memory[8057] = 32'd216;
     memory[8058] = 32'd183;
     memory[8059] = 32'd134;
     memory[8060] = 32'd31;
     memory[8061] = 32'd186;
     memory[8062] = 32'd235;
     memory[8063] = 32'd166;
     memory[8064] = 32'd54;
     memory[8065] = 32'd9;
     memory[8066] = 32'd163;
     memory[8067] = 32'd100;
     memory[8068] = 32'd128;
     memory[8069] = 32'd250;
     memory[8070] = 32'd221;
     memory[8071] = 32'd117;
     memory[8072] = 32'd16;
     memory[8073] = 32'd137;
     memory[8074] = 32'd194;
     memory[8075] = 32'd12;
     memory[8076] = 32'd61;
     memory[8077] = 32'd102;
     memory[8078] = 32'd129;
     memory[8079] = 32'd182;
     memory[8080] = 32'd38;
     memory[8081] = 32'd51;
     memory[8082] = 32'd17;
     memory[8083] = 32'd189;
     memory[8084] = 32'd222;
     memory[8085] = 32'd171;
     memory[8086] = 32'd229;
     memory[8087] = 32'd240;
     memory[8088] = 32'd248;
     memory[8089] = 32'd136;
     memory[8090] = 32'd151;
     memory[8091] = 32'd237;
     memory[8092] = 32'd218;
     memory[8093] = 32'd141;
     memory[8094] = 32'd52;
     memory[8095] = 32'd150;
     memory[8096] = 32'd30;
     memory[8097] = 32'd222;
     memory[8098] = 32'd9;
     memory[8099] = 32'd142;
     memory[8100] = 32'd142;
     memory[8101] = 32'd244;
     memory[8102] = 32'd113;
     memory[8103] = 32'd82;
     memory[8104] = 32'd43;
     memory[8105] = 32'd70;
     memory[8106] = 32'd170;
     memory[8107] = 32'd215;
     memory[8108] = 32'd251;
     memory[8109] = 32'd217;
     memory[8110] = 32'd101;
     memory[8111] = 32'd116;
     memory[8112] = 32'd71;
     memory[8113] = 32'd196;
     memory[8114] = 32'd166;
     memory[8115] = 32'd235;
     memory[8116] = 32'd147;
     memory[8117] = 32'd39;
     memory[8118] = 32'd138;
     memory[8119] = 32'd237;
     memory[8120] = 32'd179;
     memory[8121] = 32'd143;
     memory[8122] = 32'd241;
     memory[8123] = 32'd32;
     memory[8124] = 32'd174;
     memory[8125] = 32'd7;
     memory[8126] = 32'd17;
     memory[8127] = 32'd87;
     memory[8128] = 32'd31;
     memory[8129] = 32'd93;
     memory[8130] = 32'd219;
     memory[8131] = 32'd55;
     memory[8132] = 32'd97;
     memory[8133] = 32'd144;
     memory[8134] = 32'd99;
     memory[8135] = 32'd246;
     memory[8136] = 32'd115;
     memory[8137] = 32'd49;
     memory[8138] = 32'd92;
     memory[8139] = 32'd102;
     memory[8140] = 32'd49;
     memory[8141] = 32'd164;
     memory[8142] = 32'd7;
     memory[8143] = 32'd119;
     memory[8144] = 32'd116;
     memory[8145] = 32'd232;
     memory[8146] = 32'd22;
     memory[8147] = 32'd140;
     memory[8148] = 32'd80;
     memory[8149] = 32'd150;
     memory[8150] = 32'd5;
     memory[8151] = 32'd6;
     memory[8152] = 32'd100;
     memory[8153] = 32'd31;
     memory[8154] = 32'd146;
     memory[8155] = 32'd18;
     memory[8156] = 32'd184;
     memory[8157] = 32'd144;
     memory[8158] = 32'd83;
     memory[8159] = 32'd3;
     memory[8160] = 32'd18;
     memory[8161] = 32'd211;
     memory[8162] = 32'd121;
     memory[8163] = 32'd128;
     memory[8164] = 32'd137;
     memory[8165] = 32'd57;
     memory[8166] = 32'd56;
     memory[8167] = 32'd112;
     memory[8168] = 32'd113;
     memory[8169] = 32'd103;
     memory[8170] = 32'd154;
     memory[8171] = 32'd38;
     memory[8172] = 32'd163;
     memory[8173] = 32'd250;
     memory[8174] = 32'd226;
     memory[8175] = 32'd19;
     memory[8176] = 32'd172;
     memory[8177] = 32'd145;
     memory[8178] = 32'd118;
     memory[8179] = 32'd153;
     memory[8180] = 32'd1;
     memory[8181] = 32'd119;
     memory[8182] = 32'd173;
     memory[8183] = 32'd227;
     memory[8184] = 32'd139;
     memory[8185] = 32'd249;
     memory[8186] = 32'd210;
     memory[8187] = 32'd39;
     memory[8188] = 32'd32;
     memory[8189] = 32'd36;
     memory[8190] = 32'd59;
     memory[8191] = 32'd151;
     memory[8192] = 32'd146;
     memory[8193] = 32'd1;
     memory[8194] = 32'd1;
     memory[8195] = 32'd1;
     memory[8196] = 32'd1;
     memory[8197] = 32'd1;
     memory[8198] = 32'd0;
     memory[8199] = 32'd0;
     memory[8200] = 32'd1;
     memory[8201] = 32'd1;
     memory[8202] = 32'd1;
     memory[8203] = 32'd0;
     memory[8204] = 32'd1;
     memory[8205] = 32'd0;
     memory[8206] = 32'd0;
     memory[8207] = 32'd1;
     memory[8208] = 32'd0;
     memory[8209] = 32'd1;
     memory[8210] = 32'd1;
     memory[8211] = 32'd1;
     memory[8212] = 32'd1;
     memory[8213] = 32'd0;
     memory[8214] = 32'd0;
     memory[8215] = 32'd1;
     memory[8216] = 32'd1;
     memory[8217] = 32'd1;
     memory[8218] = 32'd0;
     memory[8219] = 32'd1;
     memory[8220] = 32'd1;
     memory[8221] = 32'd0;
     memory[8222] = 32'd1;
     memory[8223] = 32'd0;
     memory[8224] = 32'd0;
     memory[8225] = 32'd0;
     memory[8226] = 32'd1;
     memory[8227] = 32'd1;
     memory[8228] = 32'd0;
     memory[8229] = 32'd0;
     memory[8230] = 32'd1;
     memory[8231] = 32'd0;
     memory[8232] = 32'd0;
     memory[8233] = 32'd1;
     memory[8234] = 32'd1;
     memory[8235] = 32'd0;
     memory[8236] = 32'd0;
     memory[8237] = 32'd1;
     memory[8238] = 32'd0;
     memory[8239] = 32'd1;
     memory[8240] = 32'd0;
     memory[8241] = 32'd1;
     memory[8242] = 32'd1;
     memory[8243] = 32'd1;
     memory[8244] = 32'd1;
     memory[8245] = 32'd0;
     memory[8246] = 32'd1;
     memory[8247] = 32'd1;
     memory[8248] = 32'd0;
     memory[8249] = 32'd1;
     memory[8250] = 32'd1;
     memory[8251] = 32'd1;
     memory[8252] = 32'd0;
     memory[8253] = 32'd1;
     memory[8254] = 32'd0;
     memory[8255] = 32'd0;
     memory[8256] = 32'd0;
     memory[8257] = 32'd0;
     memory[8258] = 32'd1;
     memory[8259] = 32'd0;
     memory[8260] = 32'd0;
     memory[8261] = 32'd1;
     memory[8262] = 32'd0;
     memory[8263] = 32'd1;
     memory[8264] = 32'd0;
     memory[8265] = 32'd1;
     memory[8266] = 32'd0;
     memory[8267] = 32'd0;
     memory[8268] = 32'd0;
     memory[8269] = 32'd0;
     memory[8270] = 32'd0;
     memory[8271] = 32'd0;
     memory[8272] = 32'd0;
     memory[8273] = 32'd1;
     memory[8274] = 32'd0;
     memory[8275] = 32'd1;
     memory[8276] = 32'd1;
     memory[8277] = 32'd0;
     memory[8278] = 32'd0;
     memory[8279] = 32'd0;
     memory[8280] = 32'd1;
     memory[8281] = 32'd1;
     memory[8282] = 32'd0;
     memory[8283] = 32'd1;
     memory[8284] = 32'd1;
     memory[8285] = 32'd1;
     memory[8286] = 32'd0;
     memory[8287] = 32'd1;
     memory[8288] = 32'd1;
     memory[8289] = 32'd0;
     memory[8290] = 32'd0;
     memory[8291] = 32'd1;
     memory[8292] = 32'd0;
     memory[8293] = 32'd1;
     memory[8294] = 32'd0;
     memory[8295] = 32'd0;
     memory[8296] = 32'd0;
     memory[8297] = 32'd1;
     memory[8298] = 32'd0;
     memory[8299] = 32'd1;
     memory[8300] = 32'd1;
     memory[8301] = 32'd0;
     memory[8302] = 32'd1;
     memory[8303] = 32'd1;
     memory[8304] = 32'd0;
     memory[8305] = 32'd0;
     memory[8306] = 32'd1;
     memory[8307] = 32'd1;
     memory[8308] = 32'd0;
     memory[8309] = 32'd1;
     memory[8310] = 32'd1;
     memory[8311] = 32'd1;
     memory[8312] = 32'd0;
     memory[8313] = 32'd1;
     memory[8314] = 32'd1;
     memory[8315] = 32'd0;
     memory[8316] = 32'd1;
     memory[8317] = 32'd0;
     memory[8318] = 32'd1;
     memory[8319] = 32'd1;
     memory[8320] = 32'd1;
     memory[8321] = 32'd0;
     memory[8322] = 32'd1;
     memory[8323] = 32'd1;
     memory[8324] = 32'd1;
     memory[8325] = 32'd0;
     memory[8326] = 32'd1;
     memory[8327] = 32'd1;
     memory[8328] = 32'd1;
     memory[8329] = 32'd1;
     memory[8330] = 32'd0;
     memory[8331] = 32'd0;
     memory[8332] = 32'd0;
     memory[8333] = 32'd1;
     memory[8334] = 32'd0;
     memory[8335] = 32'd1;
     memory[8336] = 32'd1;
     memory[8337] = 32'd0;
     memory[8338] = 32'd1;
     memory[8339] = 32'd0;
     memory[8340] = 32'd1;
     memory[8341] = 32'd1;
     memory[8342] = 32'd0;
     memory[8343] = 32'd1;
     memory[8344] = 32'd0;
     memory[8345] = 32'd1;
     memory[8346] = 32'd0;
     memory[8347] = 32'd1;
     memory[8348] = 32'd0;
     memory[8349] = 32'd0;
     memory[8350] = 32'd0;
     memory[8351] = 32'd0;
     memory[8352] = 32'd1;
     memory[8353] = 32'd1;
     memory[8354] = 32'd1;
     memory[8355] = 32'd1;
     memory[8356] = 32'd1;
     memory[8357] = 32'd0;
     memory[8358] = 32'd0;
     memory[8359] = 32'd0;
     memory[8360] = 32'd1;
     memory[8361] = 32'd1;
     memory[8362] = 32'd0;
     memory[8363] = 32'd1;
     memory[8364] = 32'd0;
     memory[8365] = 32'd1;
     memory[8366] = 32'd0;
     memory[8367] = 32'd0;
     memory[8368] = 32'd0;
     memory[8369] = 32'd0;
     memory[8370] = 32'd1;
     memory[8371] = 32'd1;
     memory[8372] = 32'd1;
     memory[8373] = 32'd1;
     memory[8374] = 32'd0;
     memory[8375] = 32'd1;
     memory[8376] = 32'd1;
     memory[8377] = 32'd1;
     memory[8378] = 32'd1;
     memory[8379] = 32'd0;
     memory[8380] = 32'd1;
     memory[8381] = 32'd0;
     memory[8382] = 32'd1;
     memory[8383] = 32'd1;
     memory[8384] = 32'd0;
     memory[8385] = 32'd1;
     memory[8386] = 32'd0;
     memory[8387] = 32'd0;
     memory[8388] = 32'd1;
     memory[8389] = 32'd1;
     memory[8390] = 32'd1;
     memory[8391] = 32'd1;
     memory[8392] = 32'd1;
     memory[8393] = 32'd0;
     memory[8394] = 32'd0;
     memory[8395] = 32'd0;
     memory[8396] = 32'd0;
     memory[8397] = 32'd0;
     memory[8398] = 32'd0;
     memory[8399] = 32'd0;
     memory[8400] = 32'd0;
     memory[8401] = 32'd0;
     memory[8402] = 32'd0;
     memory[8403] = 32'd0;
     memory[8404] = 32'd0;
     memory[8405] = 32'd0;
     memory[8406] = 32'd0;
     memory[8407] = 32'd0;
     memory[8408] = 32'd0;
     memory[8409] = 32'd0;
     memory[8410] = 32'd1;
     memory[8411] = 32'd0;
     memory[8412] = 32'd1;
     memory[8413] = 32'd1;
     memory[8414] = 32'd0;
     memory[8415] = 32'd0;
     memory[8416] = 32'd0;
     memory[8417] = 32'd0;
     memory[8418] = 32'd1;
     memory[8419] = 32'd1;
     memory[8420] = 32'd1;
     memory[8421] = 32'd0;
     memory[8422] = 32'd1;
     memory[8423] = 32'd1;
     memory[8424] = 32'd1;
     memory[8425] = 32'd0;
     memory[8426] = 32'd1;
     memory[8427] = 32'd0;
     memory[8428] = 32'd0;
     memory[8429] = 32'd1;
     memory[8430] = 32'd0;
     memory[8431] = 32'd1;
     memory[8432] = 32'd1;
     memory[8433] = 32'd0;
     memory[8434] = 32'd1;
     memory[8435] = 32'd1;
     memory[8436] = 32'd1;
     memory[8437] = 32'd0;
     memory[8438] = 32'd0;
     memory[8439] = 32'd1;
     memory[8440] = 32'd0;
     memory[8441] = 32'd1;
     memory[8442] = 32'd1;
     memory[8443] = 32'd1;
     memory[8444] = 32'd1;
     memory[8445] = 32'd1;
     memory[8446] = 32'd1;
     memory[8447] = 32'd0;
     memory[8448] = 32'd0;
     memory[8449] = 32'd1;
     memory[8450] = 32'd1;
     memory[8451] = 32'd1;
     memory[8452] = 32'd1;
     memory[8453] = 32'd1;
     memory[8454] = 32'd1;
     memory[8455] = 32'd0;
     memory[8456] = 32'd0;
     memory[8457] = 32'd1;
     memory[8458] = 32'd0;
     memory[8459] = 32'd0;
     memory[8460] = 32'd1;
     memory[8461] = 32'd0;
     memory[8462] = 32'd0;
     memory[8463] = 32'd1;
     memory[8464] = 32'd1;
     memory[8465] = 32'd1;
     memory[8466] = 32'd0;
     memory[8467] = 32'd1;
     memory[8468] = 32'd0;
     memory[8469] = 32'd0;
     memory[8470] = 32'd0;
     memory[8471] = 32'd1;
     memory[8472] = 32'd0;
     memory[8473] = 32'd1;
     memory[8474] = 32'd1;
     memory[8475] = 32'd0;
     memory[8476] = 32'd1;
     memory[8477] = 32'd1;
     memory[8478] = 32'd1;
     memory[8479] = 32'd0;
     memory[8480] = 32'd1;
     memory[8481] = 32'd0;
     memory[8482] = 32'd1;
     memory[8483] = 32'd0;
     memory[8484] = 32'd1;
     memory[8485] = 32'd1;
     memory[8486] = 32'd0;
     memory[8487] = 32'd1;
     memory[8488] = 32'd1;
     memory[8489] = 32'd1;
     memory[8490] = 32'd1;
     memory[8491] = 32'd1;
     memory[8492] = 32'd0;
     memory[8493] = 32'd0;
     memory[8494] = 32'd0;
     memory[8495] = 32'd0;
     memory[8496] = 32'd1;
     memory[8497] = 32'd1;
     memory[8498] = 32'd0;
     memory[8499] = 32'd0;
     memory[8500] = 32'd0;
     memory[8501] = 32'd0;
     memory[8502] = 32'd0;
     memory[8503] = 32'd0;
     memory[8504] = 32'd1;
     memory[8505] = 32'd0;
     memory[8506] = 32'd0;
     memory[8507] = 32'd1;
     memory[8508] = 32'd0;
     memory[8509] = 32'd0;
     memory[8510] = 32'd1;
     memory[8511] = 32'd0;
     memory[8512] = 32'd0;
     memory[8513] = 32'd0;
     memory[8514] = 32'd0;
     memory[8515] = 32'd1;
     memory[8516] = 32'd1;
     memory[8517] = 32'd0;
     memory[8518] = 32'd1;
     memory[8519] = 32'd0;
     memory[8520] = 32'd0;
     memory[8521] = 32'd1;
     memory[8522] = 32'd0;
     memory[8523] = 32'd1;
     memory[8524] = 32'd1;
     memory[8525] = 32'd0;
     memory[8526] = 32'd0;
     memory[8527] = 32'd1;
     memory[8528] = 32'd0;
     memory[8529] = 32'd0;
     memory[8530] = 32'd1;
     memory[8531] = 32'd1;
     memory[8532] = 32'd0;
     memory[8533] = 32'd1;
     memory[8534] = 32'd0;
     memory[8535] = 32'd0;
     memory[8536] = 32'd1;
     memory[8537] = 32'd1;
     memory[8538] = 32'd0;
     memory[8539] = 32'd0;
     memory[8540] = 32'd0;
     memory[8541] = 32'd1;
     memory[8542] = 32'd0;
     memory[8543] = 32'd0;
     memory[8544] = 32'd1;
     memory[8545] = 32'd1;
     memory[8546] = 32'd1;
     memory[8547] = 32'd0;
     memory[8548] = 32'd0;
     memory[8549] = 32'd1;
     memory[8550] = 32'd1;
     memory[8551] = 32'd0;
     memory[8552] = 32'd0;
     memory[8553] = 32'd1;
     memory[8554] = 32'd1;
     memory[8555] = 32'd0;
     memory[8556] = 32'd0;
     memory[8557] = 32'd0;
     memory[8558] = 32'd1;
     memory[8559] = 32'd0;
     memory[8560] = 32'd1;
     memory[8561] = 32'd0;
     memory[8562] = 32'd1;
     memory[8563] = 32'd0;
     memory[8564] = 32'd1;
     memory[8565] = 32'd0;
     memory[8566] = 32'd0;
     memory[8567] = 32'd0;
     memory[8568] = 32'd1;
     memory[8569] = 32'd0;
     memory[8570] = 32'd0;
     memory[8571] = 32'd0;
     memory[8572] = 32'd1;
     memory[8573] = 32'd1;
     memory[8574] = 32'd1;
     memory[8575] = 32'd1;
     memory[8576] = 32'd1;
     memory[8577] = 32'd1;
     memory[8578] = 32'd1;
     memory[8579] = 32'd0;
     memory[8580] = 32'd1;
     memory[8581] = 32'd0;
     memory[8582] = 32'd0;
     memory[8583] = 32'd1;
     memory[8584] = 32'd1;
     memory[8585] = 32'd1;
     memory[8586] = 32'd0;
     memory[8587] = 32'd0;
     memory[8588] = 32'd0;
     memory[8589] = 32'd1;
     memory[8590] = 32'd1;
     memory[8591] = 32'd1;
     memory[8592] = 32'd1;
     memory[8593] = 32'd0;
     memory[8594] = 32'd1;
     memory[8595] = 32'd0;
     memory[8596] = 32'd1;
     memory[8597] = 32'd0;
     memory[8598] = 32'd0;
     memory[8599] = 32'd1;
     memory[8600] = 32'd0;
     memory[8601] = 32'd0;
     memory[8602] = 32'd0;
     memory[8603] = 32'd0;
     memory[8604] = 32'd0;
     memory[8605] = 32'd1;
     memory[8606] = 32'd0;
     memory[8607] = 32'd0;
     memory[8608] = 32'd1;
     memory[8609] = 32'd1;
     memory[8610] = 32'd1;
     memory[8611] = 32'd0;
     memory[8612] = 32'd1;
     memory[8613] = 32'd1;
     memory[8614] = 32'd0;
     memory[8615] = 32'd0;
     memory[8616] = 32'd1;
     memory[8617] = 32'd0;
     memory[8618] = 32'd0;
     memory[8619] = 32'd1;
     memory[8620] = 32'd0;
     memory[8621] = 32'd1;
     memory[8622] = 32'd1;
     memory[8623] = 32'd0;
     memory[8624] = 32'd0;
     memory[8625] = 32'd0;
     memory[8626] = 32'd0;
     memory[8627] = 32'd0;
     memory[8628] = 32'd0;
     memory[8629] = 32'd1;
     memory[8630] = 32'd1;
     memory[8631] = 32'd0;
     memory[8632] = 32'd1;
     memory[8633] = 32'd1;
     memory[8634] = 32'd1;
     memory[8635] = 32'd1;
     memory[8636] = 32'd0;
     memory[8637] = 32'd0;
     memory[8638] = 32'd1;
     memory[8639] = 32'd0;
     memory[8640] = 32'd0;
     memory[8641] = 32'd0;
     memory[8642] = 32'd0;
     memory[8643] = 32'd0;
     memory[8644] = 32'd1;
     memory[8645] = 32'd1;
     memory[8646] = 32'd0;
     memory[8647] = 32'd1;
     memory[8648] = 32'd1;
     memory[8649] = 32'd0;
     memory[8650] = 32'd0;
     memory[8651] = 32'd1;
     memory[8652] = 32'd1;
     memory[8653] = 32'd0;
     memory[8654] = 32'd0;
     memory[8655] = 32'd0;
     memory[8656] = 32'd0;
     memory[8657] = 32'd0;
     memory[8658] = 32'd1;
     memory[8659] = 32'd0;
     memory[8660] = 32'd0;
     memory[8661] = 32'd0;
     memory[8662] = 32'd0;
     memory[8663] = 32'd1;
     memory[8664] = 32'd1;
     memory[8665] = 32'd0;
     memory[8666] = 32'd1;
     memory[8667] = 32'd1;
     memory[8668] = 32'd1;
     memory[8669] = 32'd0;
     memory[8670] = 32'd0;
     memory[8671] = 32'd0;
     memory[8672] = 32'd0;
     memory[8673] = 32'd1;
     memory[8674] = 32'd0;
     memory[8675] = 32'd1;
     memory[8676] = 32'd1;
     memory[8677] = 32'd1;
     memory[8678] = 32'd1;
     memory[8679] = 32'd0;
     memory[8680] = 32'd1;
     memory[8681] = 32'd0;
     memory[8682] = 32'd1;
     memory[8683] = 32'd1;
     memory[8684] = 32'd1;
     memory[8685] = 32'd1;
     memory[8686] = 32'd0;
     memory[8687] = 32'd1;
     memory[8688] = 32'd1;
     memory[8689] = 32'd1;
     memory[8690] = 32'd1;
     memory[8691] = 32'd1;
     memory[8692] = 32'd0;
     memory[8693] = 32'd1;
     memory[8694] = 32'd0;
     memory[8695] = 32'd0;
     memory[8696] = 32'd0;
     memory[8697] = 32'd0;
     memory[8698] = 32'd0;
     memory[8699] = 32'd1;
     memory[8700] = 32'd0;
     memory[8701] = 32'd1;
     memory[8702] = 32'd0;
     memory[8703] = 32'd1;
     memory[8704] = 32'd1;
     memory[8705] = 32'd0;
     memory[8706] = 32'd1;
     memory[8707] = 32'd1;
     memory[8708] = 32'd0;
     memory[8709] = 32'd1;
     memory[8710] = 32'd0;
     memory[8711] = 32'd0;
     memory[8712] = 32'd0;
     memory[8713] = 32'd1;
     memory[8714] = 32'd0;
     memory[8715] = 32'd1;
     memory[8716] = 32'd1;
     memory[8717] = 32'd1;
     memory[8718] = 32'd1;
     memory[8719] = 32'd1;
     memory[8720] = 32'd0;
     memory[8721] = 32'd1;
     memory[8722] = 32'd1;
     memory[8723] = 32'd1;
     memory[8724] = 32'd1;
     memory[8725] = 32'd0;
     memory[8726] = 32'd0;
     memory[8727] = 32'd1;
     memory[8728] = 32'd0;
     memory[8729] = 32'd1;
     memory[8730] = 32'd0;
     memory[8731] = 32'd1;
     memory[8732] = 32'd0;
     memory[8733] = 32'd1;
     memory[8734] = 32'd1;
     memory[8735] = 32'd0;
     memory[8736] = 32'd0;
     memory[8737] = 32'd0;
     memory[8738] = 32'd0;
     memory[8739] = 32'd0;
     memory[8740] = 32'd0;
     memory[8741] = 32'd1;
     memory[8742] = 32'd0;
     memory[8743] = 32'd0;
     memory[8744] = 32'd0;
     memory[8745] = 32'd0;
     memory[8746] = 32'd0;
     memory[8747] = 32'd1;
     memory[8748] = 32'd0;
     memory[8749] = 32'd1;
     memory[8750] = 32'd1;
     memory[8751] = 32'd0;
     memory[8752] = 32'd0;
     memory[8753] = 32'd0;
     memory[8754] = 32'd1;
     memory[8755] = 32'd0;
     memory[8756] = 32'd1;
     memory[8757] = 32'd1;
     memory[8758] = 32'd0;
     memory[8759] = 32'd0;
     memory[8760] = 32'd1;
     memory[8761] = 32'd1;
     memory[8762] = 32'd1;
     memory[8763] = 32'd1;
     memory[8764] = 32'd0;
     memory[8765] = 32'd0;
     memory[8766] = 32'd0;
     memory[8767] = 32'd1;
     memory[8768] = 32'd0;
     memory[8769] = 32'd1;
     memory[8770] = 32'd0;
     memory[8771] = 32'd0;
     memory[8772] = 32'd1;
     memory[8773] = 32'd1;
     memory[8774] = 32'd1;
     memory[8775] = 32'd1;
     memory[8776] = 32'd0;
     memory[8777] = 32'd1;
     memory[8778] = 32'd0;
     memory[8779] = 32'd0;
     memory[8780] = 32'd0;
     memory[8781] = 32'd0;
     memory[8782] = 32'd1;
     memory[8783] = 32'd0;
     memory[8784] = 32'd0;
     memory[8785] = 32'd1;
     memory[8786] = 32'd1;
     memory[8787] = 32'd0;
     memory[8788] = 32'd0;
     memory[8789] = 32'd1;
     memory[8790] = 32'd1;
     memory[8791] = 32'd1;
     memory[8792] = 32'd1;
     memory[8793] = 32'd1;
     memory[8794] = 32'd1;
     memory[8795] = 32'd1;
     memory[8796] = 32'd0;
     memory[8797] = 32'd1;
     memory[8798] = 32'd0;
     memory[8799] = 32'd1;
     memory[8800] = 32'd1;
     memory[8801] = 32'd1;
     memory[8802] = 32'd1;
     memory[8803] = 32'd0;
     memory[8804] = 32'd0;
     memory[8805] = 32'd0;
     memory[8806] = 32'd0;
     memory[8807] = 32'd0;
     memory[8808] = 32'd1;
     memory[8809] = 32'd0;
     memory[8810] = 32'd1;
     memory[8811] = 32'd1;
     memory[8812] = 32'd1;
     memory[8813] = 32'd1;
     memory[8814] = 32'd0;
     memory[8815] = 32'd1;
     memory[8816] = 32'd0;
     memory[8817] = 32'd0;
     memory[8818] = 32'd1;
     memory[8819] = 32'd0;
     memory[8820] = 32'd0;
     memory[8821] = 32'd0;
     memory[8822] = 32'd0;
     memory[8823] = 32'd0;
     memory[8824] = 32'd1;
     memory[8825] = 32'd0;
     memory[8826] = 32'd1;
     memory[8827] = 32'd1;
     memory[8828] = 32'd1;
     memory[8829] = 32'd1;
     memory[8830] = 32'd0;
     memory[8831] = 32'd1;
     memory[8832] = 32'd1;
     memory[8833] = 32'd0;
     memory[8834] = 32'd0;
     memory[8835] = 32'd1;
     memory[8836] = 32'd0;
     memory[8837] = 32'd1;
     memory[8838] = 32'd1;
     memory[8839] = 32'd0;
     memory[8840] = 32'd1;
     memory[8841] = 32'd0;
     memory[8842] = 32'd0;
     memory[8843] = 32'd1;
     memory[8844] = 32'd0;
     memory[8845] = 32'd1;
     memory[8846] = 32'd1;
     memory[8847] = 32'd0;
     memory[8848] = 32'd1;
     memory[8849] = 32'd0;
     memory[8850] = 32'd0;
     memory[8851] = 32'd0;
     memory[8852] = 32'd0;
     memory[8853] = 32'd1;
     memory[8854] = 32'd0;
     memory[8855] = 32'd1;
     memory[8856] = 32'd0;
     memory[8857] = 32'd0;
     memory[8858] = 32'd1;
     memory[8859] = 32'd0;
     memory[8860] = 32'd1;
     memory[8861] = 32'd0;
     memory[8862] = 32'd0;
     memory[8863] = 32'd0;
     memory[8864] = 32'd0;
     memory[8865] = 32'd0;
     memory[8866] = 32'd0;
     memory[8867] = 32'd0;
     memory[8868] = 32'd1;
     memory[8869] = 32'd1;
     memory[8870] = 32'd0;
     memory[8871] = 32'd0;
     memory[8872] = 32'd1;
     memory[8873] = 32'd1;
     memory[8874] = 32'd1;
     memory[8875] = 32'd0;
     memory[8876] = 32'd1;
     memory[8877] = 32'd0;
     memory[8878] = 32'd1;
     memory[8879] = 32'd1;
     memory[8880] = 32'd0;
     memory[8881] = 32'd1;
     memory[8882] = 32'd0;
     memory[8883] = 32'd1;
     memory[8884] = 32'd0;
     memory[8885] = 32'd0;
     memory[8886] = 32'd1;
     memory[8887] = 32'd1;
     memory[8888] = 32'd0;
     memory[8889] = 32'd1;
     memory[8890] = 32'd0;
     memory[8891] = 32'd1;
     memory[8892] = 32'd1;
     memory[8893] = 32'd0;
     memory[8894] = 32'd0;
     memory[8895] = 32'd1;
     memory[8896] = 32'd1;
     memory[8897] = 32'd0;
     memory[8898] = 32'd0;
     memory[8899] = 32'd1;
     memory[8900] = 32'd0;
     memory[8901] = 32'd1;
     memory[8902] = 32'd1;
     memory[8903] = 32'd0;
     memory[8904] = 32'd1;
     memory[8905] = 32'd0;
     memory[8906] = 32'd0;
     memory[8907] = 32'd0;
     memory[8908] = 32'd1;
     memory[8909] = 32'd1;
     memory[8910] = 32'd0;
     memory[8911] = 32'd1;
     memory[8912] = 32'd0;
     memory[8913] = 32'd0;
     memory[8914] = 32'd0;
     memory[8915] = 32'd1;
     memory[8916] = 32'd0;
     memory[8917] = 32'd0;
     memory[8918] = 32'd1;
     memory[8919] = 32'd1;
     memory[8920] = 32'd1;
     memory[8921] = 32'd0;
     memory[8922] = 32'd1;
     memory[8923] = 32'd1;
     memory[8924] = 32'd0;
     memory[8925] = 32'd0;
     memory[8926] = 32'd1;
     memory[8927] = 32'd0;
     memory[8928] = 32'd1;
     memory[8929] = 32'd0;
     memory[8930] = 32'd0;
     memory[8931] = 32'd1;
     memory[8932] = 32'd1;
     memory[8933] = 32'd0;
     memory[8934] = 32'd0;
     memory[8935] = 32'd1;
     memory[8936] = 32'd1;
     memory[8937] = 32'd0;
     memory[8938] = 32'd0;
     memory[8939] = 32'd0;
     memory[8940] = 32'd1;
     memory[8941] = 32'd1;
     memory[8942] = 32'd1;
     memory[8943] = 32'd0;
     memory[8944] = 32'd1;
     memory[8945] = 32'd0;
     memory[8946] = 32'd1;
     memory[8947] = 32'd1;
     memory[8948] = 32'd1;
     memory[8949] = 32'd1;
     memory[8950] = 32'd0;
     memory[8951] = 32'd0;
     memory[8952] = 32'd0;
     memory[8953] = 32'd0;
     memory[8954] = 32'd0;
     memory[8955] = 32'd0;
     memory[8956] = 32'd0;
     memory[8957] = 32'd1;
     memory[8958] = 32'd1;
     memory[8959] = 32'd0;
     memory[8960] = 32'd0;
     memory[8961] = 32'd0;
     memory[8962] = 32'd1;
     memory[8963] = 32'd0;
     memory[8964] = 32'd0;
     memory[8965] = 32'd0;
     memory[8966] = 32'd1;
     memory[8967] = 32'd1;
     memory[8968] = 32'd0;
     memory[8969] = 32'd1;
     memory[8970] = 32'd0;
     memory[8971] = 32'd1;
     memory[8972] = 32'd1;
     memory[8973] = 32'd1;
     memory[8974] = 32'd1;
     memory[8975] = 32'd1;
     memory[8976] = 32'd0;
     memory[8977] = 32'd1;
     memory[8978] = 32'd1;
     memory[8979] = 32'd1;
     memory[8980] = 32'd1;
     memory[8981] = 32'd0;
     memory[8982] = 32'd0;
     memory[8983] = 32'd0;
     memory[8984] = 32'd0;
     memory[8985] = 32'd0;
     memory[8986] = 32'd0;
     memory[8987] = 32'd0;
     memory[8988] = 32'd0;
     memory[8989] = 32'd0;
     memory[8990] = 32'd1;
     memory[8991] = 32'd0;
     memory[8992] = 32'd1;
     memory[8993] = 32'd1;
     memory[8994] = 32'd0;
     memory[8995] = 32'd1;
     memory[8996] = 32'd1;
     memory[8997] = 32'd1;
     memory[8998] = 32'd1;
     memory[8999] = 32'd1;
     memory[9000] = 32'd0;
     memory[9001] = 32'd0;
     memory[9002] = 32'd0;
     memory[9003] = 32'd1;
     memory[9004] = 32'd0;
     memory[9005] = 32'd0;
     memory[9006] = 32'd1;
     memory[9007] = 32'd1;
     memory[9008] = 32'd1;
     memory[9009] = 32'd0;
     memory[9010] = 32'd1;
     memory[9011] = 32'd0;
     memory[9012] = 32'd1;
     memory[9013] = 32'd1;
     memory[9014] = 32'd1;
     memory[9015] = 32'd1;
     memory[9016] = 32'd0;
     memory[9017] = 32'd1;
     memory[9018] = 32'd1;
     memory[9019] = 32'd1;
     memory[9020] = 32'd1;
     memory[9021] = 32'd1;
     memory[9022] = 32'd0;
     memory[9023] = 32'd0;
     memory[9024] = 32'd0;
     memory[9025] = 32'd0;
     memory[9026] = 32'd0;
     memory[9027] = 32'd1;
     memory[9028] = 32'd0;
     memory[9029] = 32'd1;
     memory[9030] = 32'd1;
     memory[9031] = 32'd1;
     memory[9032] = 32'd0;
     memory[9033] = 32'd0;
     memory[9034] = 32'd0;
     memory[9035] = 32'd0;
     memory[9036] = 32'd0;
     memory[9037] = 32'd1;
     memory[9038] = 32'd1;
     memory[9039] = 32'd1;
     memory[9040] = 32'd0;
     memory[9041] = 32'd0;
     memory[9042] = 32'd1;
     memory[9043] = 32'd0;
     memory[9044] = 32'd1;
     memory[9045] = 32'd0;
     memory[9046] = 32'd1;
     memory[9047] = 32'd0;
     memory[9048] = 32'd1;
     memory[9049] = 32'd0;
     memory[9050] = 32'd0;
     memory[9051] = 32'd0;
     memory[9052] = 32'd1;
     memory[9053] = 32'd1;
     memory[9054] = 32'd1;
     memory[9055] = 32'd0;
     memory[9056] = 32'd0;
     memory[9057] = 32'd0;
     memory[9058] = 32'd0;
     memory[9059] = 32'd1;
     memory[9060] = 32'd1;
     memory[9061] = 32'd0;
     memory[9062] = 32'd1;
     memory[9063] = 32'd1;
     memory[9064] = 32'd1;
     memory[9065] = 32'd0;
     memory[9066] = 32'd1;
     memory[9067] = 32'd1;
     memory[9068] = 32'd0;
     memory[9069] = 32'd1;
     memory[9070] = 32'd0;
     memory[9071] = 32'd1;
     memory[9072] = 32'd1;
     memory[9073] = 32'd1;
     memory[9074] = 32'd1;
     memory[9075] = 32'd0;
     memory[9076] = 32'd1;
     memory[9077] = 32'd0;
     memory[9078] = 32'd1;
     memory[9079] = 32'd0;
     memory[9080] = 32'd0;
     memory[9081] = 32'd0;
     memory[9082] = 32'd0;
     memory[9083] = 32'd1;
     memory[9084] = 32'd0;
     memory[9085] = 32'd0;
     memory[9086] = 32'd1;
     memory[9087] = 32'd1;
     memory[9088] = 32'd1;
     memory[9089] = 32'd0;
     memory[9090] = 32'd1;
     memory[9091] = 32'd0;
     memory[9092] = 32'd0;
     memory[9093] = 32'd0;
     memory[9094] = 32'd1;
     memory[9095] = 32'd1;
     memory[9096] = 32'd0;
     memory[9097] = 32'd1;
     memory[9098] = 32'd1;
     memory[9099] = 32'd1;
     memory[9100] = 32'd0;
     memory[9101] = 32'd1;
     memory[9102] = 32'd0;
     memory[9103] = 32'd0;
     memory[9104] = 32'd1;
     memory[9105] = 32'd1;
     memory[9106] = 32'd1;
     memory[9107] = 32'd1;
     memory[9108] = 32'd1;
     memory[9109] = 32'd1;
     memory[9110] = 32'd1;
     memory[9111] = 32'd0;
     memory[9112] = 32'd1;
     memory[9113] = 32'd1;
     memory[9114] = 32'd1;
     memory[9115] = 32'd0;
     memory[9116] = 32'd1;
     memory[9117] = 32'd1;
     memory[9118] = 32'd0;
     memory[9119] = 32'd0;
     memory[9120] = 32'd0;
     memory[9121] = 32'd1;
     memory[9122] = 32'd1;
     memory[9123] = 32'd0;
     memory[9124] = 32'd0;
     memory[9125] = 32'd1;
     memory[9126] = 32'd1;
     memory[9127] = 32'd1;
     memory[9128] = 32'd1;
     memory[9129] = 32'd1;
     memory[9130] = 32'd1;
     memory[9131] = 32'd0;
     memory[9132] = 32'd1;
     memory[9133] = 32'd0;
     memory[9134] = 32'd1;
     memory[9135] = 32'd1;
     memory[9136] = 32'd1;
     memory[9137] = 32'd1;
     memory[9138] = 32'd1;
     memory[9139] = 32'd1;
     memory[9140] = 32'd0;
     memory[9141] = 32'd0;
     memory[9142] = 32'd1;
     memory[9143] = 32'd1;
     memory[9144] = 32'd0;
     memory[9145] = 32'd1;
     memory[9146] = 32'd1;
     memory[9147] = 32'd1;
     memory[9148] = 32'd0;
     memory[9149] = 32'd1;
     memory[9150] = 32'd0;
     memory[9151] = 32'd1;
     memory[9152] = 32'd1;
     memory[9153] = 32'd0;
     memory[9154] = 32'd1;
     memory[9155] = 32'd1;
     memory[9156] = 32'd1;
     memory[9157] = 32'd0;
     memory[9158] = 32'd0;
     memory[9159] = 32'd1;
     memory[9160] = 32'd1;
     memory[9161] = 32'd1;
     memory[9162] = 32'd0;
     memory[9163] = 32'd1;
     memory[9164] = 32'd1;
     memory[9165] = 32'd0;
     memory[9166] = 32'd1;
     memory[9167] = 32'd0;
     memory[9168] = 32'd0;
     memory[9169] = 32'd0;
     memory[9170] = 32'd0;
     memory[9171] = 32'd1;
     memory[9172] = 32'd1;
     memory[9173] = 32'd1;
     memory[9174] = 32'd1;
     memory[9175] = 32'd0;
     memory[9176] = 32'd0;
     memory[9177] = 32'd1;
     memory[9178] = 32'd1;
     memory[9179] = 32'd0;
     memory[9180] = 32'd0;
     memory[9181] = 32'd1;
     memory[9182] = 32'd0;
     memory[9183] = 32'd1;
     memory[9184] = 32'd1;
     memory[9185] = 32'd0;
     memory[9186] = 32'd1;
     memory[9187] = 32'd0;
     memory[9188] = 32'd1;
     memory[9189] = 32'd1;
     memory[9190] = 32'd1;
     memory[9191] = 32'd1;
     memory[9192] = 32'd0;
     memory[9193] = 32'd0;
     memory[9194] = 32'd0;
     memory[9195] = 32'd1;
     memory[9196] = 32'd0;
     memory[9197] = 32'd0;
     memory[9198] = 32'd1;
     memory[9199] = 32'd0;
     memory[9200] = 32'd1;
     memory[9201] = 32'd1;
     memory[9202] = 32'd0;
     memory[9203] = 32'd1;
     memory[9204] = 32'd1;
     memory[9205] = 32'd1;
     memory[9206] = 32'd1;
     memory[9207] = 32'd1;
     memory[9208] = 32'd1;
     memory[9209] = 32'd1;
     memory[9210] = 32'd1;
     memory[9211] = 32'd1;
     memory[9212] = 32'd0;
     memory[9213] = 32'd1;
     memory[9214] = 32'd1;
     memory[9215] = 32'd1;
     memory[9216] = 32'd1;
     memory[9217] = 32'd0;
     memory[9218] = 32'd0;
     memory[9219] = 32'd1;
     memory[9220] = 32'd1;
     memory[9221] = 32'd1;
     memory[9222] = 32'd0;
     memory[9223] = 32'd0;
     memory[9224] = 32'd1;
     memory[9225] = 32'd1;
     memory[9226] = 32'd1;
     memory[9227] = 32'd0;
     memory[9228] = 32'd0;
     memory[9229] = 32'd0;
     memory[9230] = 32'd1;
     memory[9231] = 32'd0;
     memory[9232] = 32'd1;
     memory[9233] = 32'd1;
     memory[9234] = 32'd0;
     memory[9235] = 32'd1;
     memory[9236] = 32'd0;
     memory[9237] = 32'd0;
     memory[9238] = 32'd0;
     memory[9239] = 32'd1;
     memory[9240] = 32'd1;
     memory[9241] = 32'd0;
     memory[9242] = 32'd1;
     memory[9243] = 32'd1;
     memory[9244] = 32'd1;
     memory[9245] = 32'd1;
     memory[9246] = 32'd1;
     memory[9247] = 32'd0;
     memory[9248] = 32'd0;
     memory[9249] = 32'd1;
     memory[9250] = 32'd0;
     memory[9251] = 32'd0;
     memory[9252] = 32'd1;
     memory[9253] = 32'd1;
     memory[9254] = 32'd1;
     memory[9255] = 32'd1;
     memory[9256] = 32'd0;
     memory[9257] = 32'd1;
     memory[9258] = 32'd1;
     memory[9259] = 32'd0;
     memory[9260] = 32'd1;
     memory[9261] = 32'd1;
     memory[9262] = 32'd1;
     memory[9263] = 32'd0;
     memory[9264] = 32'd0;
     memory[9265] = 32'd0;
     memory[9266] = 32'd1;
     memory[9267] = 32'd1;
     memory[9268] = 32'd1;
     memory[9269] = 32'd0;
     memory[9270] = 32'd0;
     memory[9271] = 32'd0;
     memory[9272] = 32'd1;
     memory[9273] = 32'd1;
     memory[9274] = 32'd0;
     memory[9275] = 32'd1;
     memory[9276] = 32'd1;
     memory[9277] = 32'd1;
     memory[9278] = 32'd0;
     memory[9279] = 32'd0;
     memory[9280] = 32'd1;
     memory[9281] = 32'd0;
     memory[9282] = 32'd0;
     memory[9283] = 32'd1;
     memory[9284] = 32'd1;
     memory[9285] = 32'd1;
     memory[9286] = 32'd1;
     memory[9287] = 32'd1;
     memory[9288] = 32'd0;
     memory[9289] = 32'd1;
     memory[9290] = 32'd1;
     memory[9291] = 32'd1;
     memory[9292] = 32'd0;
     memory[9293] = 32'd0;
     memory[9294] = 32'd1;
     memory[9295] = 32'd1;
     memory[9296] = 32'd1;
     memory[9297] = 32'd1;
     memory[9298] = 32'd1;
     memory[9299] = 32'd0;
     memory[9300] = 32'd0;
     memory[9301] = 32'd0;
     memory[9302] = 32'd1;
     memory[9303] = 32'd1;
     memory[9304] = 32'd0;
     memory[9305] = 32'd1;
     memory[9306] = 32'd1;
     memory[9307] = 32'd1;
     memory[9308] = 32'd1;
     memory[9309] = 32'd1;
     memory[9310] = 32'd1;
     memory[9311] = 32'd1;
     memory[9312] = 32'd0;
     memory[9313] = 32'd0;
     memory[9314] = 32'd1;
     memory[9315] = 32'd0;
     memory[9316] = 32'd0;
     memory[9317] = 32'd1;
     memory[9318] = 32'd1;
     memory[9319] = 32'd1;
     memory[9320] = 32'd1;
     memory[9321] = 32'd0;
     memory[9322] = 32'd0;
     memory[9323] = 32'd1;
     memory[9324] = 32'd0;
     memory[9325] = 32'd1;
     memory[9326] = 32'd1;
     memory[9327] = 32'd0;
     memory[9328] = 32'd1;
     memory[9329] = 32'd1;
     memory[9330] = 32'd1;
     memory[9331] = 32'd0;
     memory[9332] = 32'd0;
     memory[9333] = 32'd0;
     memory[9334] = 32'd1;
     memory[9335] = 32'd0;
     memory[9336] = 32'd1;
     memory[9337] = 32'd0;
     memory[9338] = 32'd1;
     memory[9339] = 32'd1;
     memory[9340] = 32'd1;
     memory[9341] = 32'd0;
     memory[9342] = 32'd1;
     memory[9343] = 32'd0;
     memory[9344] = 32'd0;
     memory[9345] = 32'd1;
     memory[9346] = 32'd1;
     memory[9347] = 32'd0;
     memory[9348] = 32'd1;
     memory[9349] = 32'd1;
     memory[9350] = 32'd1;
     memory[9351] = 32'd0;
     memory[9352] = 32'd0;
     memory[9353] = 32'd0;
     memory[9354] = 32'd1;
     memory[9355] = 32'd0;
     memory[9356] = 32'd1;
     memory[9357] = 32'd1;
     memory[9358] = 32'd0;
     memory[9359] = 32'd1;
     memory[9360] = 32'd0;
     memory[9361] = 32'd0;
     memory[9362] = 32'd1;
     memory[9363] = 32'd1;
     memory[9364] = 32'd1;
     memory[9365] = 32'd1;
     memory[9366] = 32'd0;
     memory[9367] = 32'd1;
     memory[9368] = 32'd1;
     memory[9369] = 32'd1;
     memory[9370] = 32'd1;
     memory[9371] = 32'd1;
     memory[9372] = 32'd1;
     memory[9373] = 32'd1;
     memory[9374] = 32'd0;
     memory[9375] = 32'd0;
     memory[9376] = 32'd0;
     memory[9377] = 32'd0;
     memory[9378] = 32'd1;
     memory[9379] = 32'd0;
     memory[9380] = 32'd0;
     memory[9381] = 32'd1;
     memory[9382] = 32'd1;
     memory[9383] = 32'd1;
     memory[9384] = 32'd1;
     memory[9385] = 32'd0;
     memory[9386] = 32'd0;
     memory[9387] = 32'd0;
     memory[9388] = 32'd0;
     memory[9389] = 32'd0;
     memory[9390] = 32'd0;
     memory[9391] = 32'd1;
     memory[9392] = 32'd1;
     memory[9393] = 32'd0;
     memory[9394] = 32'd1;
     memory[9395] = 32'd1;
     memory[9396] = 32'd0;
     memory[9397] = 32'd1;
     memory[9398] = 32'd1;
     memory[9399] = 32'd1;
     memory[9400] = 32'd0;
     memory[9401] = 32'd0;
     memory[9402] = 32'd0;
     memory[9403] = 32'd1;
     memory[9404] = 32'd0;
     memory[9405] = 32'd1;
     memory[9406] = 32'd0;
     memory[9407] = 32'd0;
     memory[9408] = 32'd1;
     memory[9409] = 32'd1;
     memory[9410] = 32'd0;
     memory[9411] = 32'd1;
     memory[9412] = 32'd1;
     memory[9413] = 32'd1;
     memory[9414] = 32'd0;
     memory[9415] = 32'd1;
     memory[9416] = 32'd0;
     memory[9417] = 32'd0;
     memory[9418] = 32'd0;
     memory[9419] = 32'd1;
     memory[9420] = 32'd0;
     memory[9421] = 32'd1;
     memory[9422] = 32'd1;
     memory[9423] = 32'd1;
     memory[9424] = 32'd1;
     memory[9425] = 32'd0;
     memory[9426] = 32'd1;
     memory[9427] = 32'd1;
     memory[9428] = 32'd0;
     memory[9429] = 32'd0;
     memory[9430] = 32'd1;
     memory[9431] = 32'd1;
     memory[9432] = 32'd0;
     memory[9433] = 32'd0;
     memory[9434] = 32'd1;
     memory[9435] = 32'd0;
     memory[9436] = 32'd1;
     memory[9437] = 32'd1;
     memory[9438] = 32'd0;
     memory[9439] = 32'd0;
     memory[9440] = 32'd1;
     memory[9441] = 32'd1;
     memory[9442] = 32'd1;
     memory[9443] = 32'd1;
     memory[9444] = 32'd0;
     memory[9445] = 32'd1;
     memory[9446] = 32'd0;
     memory[9447] = 32'd1;
     memory[9448] = 32'd0;
     memory[9449] = 32'd0;
     memory[9450] = 32'd0;
     memory[9451] = 32'd0;
     memory[9452] = 32'd0;
     memory[9453] = 32'd0;
     memory[9454] = 32'd0;
     memory[9455] = 32'd1;
     memory[9456] = 32'd1;
     memory[9457] = 32'd1;
     memory[9458] = 32'd1;
     memory[9459] = 32'd1;
     memory[9460] = 32'd0;
     memory[9461] = 32'd1;
     memory[9462] = 32'd0;
     memory[9463] = 32'd0;
     memory[9464] = 32'd1;
     memory[9465] = 32'd0;
     memory[9466] = 32'd0;
     memory[9467] = 32'd0;
     memory[9468] = 32'd0;
     memory[9469] = 32'd1;
     memory[9470] = 32'd0;
     memory[9471] = 32'd0;
     memory[9472] = 32'd1;
     memory[9473] = 32'd1;
     memory[9474] = 32'd0;
     memory[9475] = 32'd1;
     memory[9476] = 32'd1;
     memory[9477] = 32'd0;
     memory[9478] = 32'd1;
     memory[9479] = 32'd0;
     memory[9480] = 32'd0;
     memory[9481] = 32'd0;
     memory[9482] = 32'd1;
     memory[9483] = 32'd0;
     memory[9484] = 32'd1;
     memory[9485] = 32'd0;
     memory[9486] = 32'd1;
     memory[9487] = 32'd0;
     memory[9488] = 32'd0;
     memory[9489] = 32'd0;
     memory[9490] = 32'd1;
     memory[9491] = 32'd1;
     memory[9492] = 32'd0;
     memory[9493] = 32'd0;
     memory[9494] = 32'd0;
     memory[9495] = 32'd0;
     memory[9496] = 32'd0;
     memory[9497] = 32'd0;
     memory[9498] = 32'd0;
     memory[9499] = 32'd0;
     memory[9500] = 32'd1;
     memory[9501] = 32'd1;
     memory[9502] = 32'd1;
     memory[9503] = 32'd1;
     memory[9504] = 32'd0;
     memory[9505] = 32'd0;
     memory[9506] = 32'd0;
     memory[9507] = 32'd0;
     memory[9508] = 32'd0;
     memory[9509] = 32'd0;
     memory[9510] = 32'd1;
     memory[9511] = 32'd0;
     memory[9512] = 32'd1;
     memory[9513] = 32'd0;
     memory[9514] = 32'd0;
     memory[9515] = 32'd1;
     memory[9516] = 32'd0;
     memory[9517] = 32'd0;
     memory[9518] = 32'd0;
     memory[9519] = 32'd0;
     memory[9520] = 32'd1;
     memory[9521] = 32'd1;
     memory[9522] = 32'd0;
     memory[9523] = 32'd1;
     memory[9524] = 32'd1;
     memory[9525] = 32'd0;
     memory[9526] = 32'd0;
     memory[9527] = 32'd1;
     memory[9528] = 32'd0;
     memory[9529] = 32'd1;
     memory[9530] = 32'd1;
     memory[9531] = 32'd1;
     memory[9532] = 32'd1;
     memory[9533] = 32'd1;
     memory[9534] = 32'd0;
     memory[9535] = 32'd0;
     memory[9536] = 32'd1;
     memory[9537] = 32'd0;
     memory[9538] = 32'd0;
     memory[9539] = 32'd0;
     memory[9540] = 32'd1;
     memory[9541] = 32'd1;
     memory[9542] = 32'd0;
     memory[9543] = 32'd0;
     memory[9544] = 32'd0;
     memory[9545] = 32'd1;
     memory[9546] = 32'd0;
     memory[9547] = 32'd1;
     memory[9548] = 32'd0;
     memory[9549] = 32'd1;
     memory[9550] = 32'd0;
     memory[9551] = 32'd1;
     memory[9552] = 32'd0;
     memory[9553] = 32'd0;
     memory[9554] = 32'd1;
     memory[9555] = 32'd0;
     memory[9556] = 32'd0;
     memory[9557] = 32'd0;
     memory[9558] = 32'd1;
     memory[9559] = 32'd1;
     memory[9560] = 32'd0;
     memory[9561] = 32'd0;
     memory[9562] = 32'd1;
     memory[9563] = 32'd1;
     memory[9564] = 32'd0;
     memory[9565] = 32'd0;
     memory[9566] = 32'd1;
     memory[9567] = 32'd1;
     memory[9568] = 32'd0;
     memory[9569] = 32'd0;
     memory[9570] = 32'd1;
     memory[9571] = 32'd1;
     memory[9572] = 32'd0;
     memory[9573] = 32'd1;
     memory[9574] = 32'd1;
     memory[9575] = 32'd1;
     memory[9576] = 32'd1;
     memory[9577] = 32'd1;
     memory[9578] = 32'd1;
     memory[9579] = 32'd1;
     memory[9580] = 32'd0;
     memory[9581] = 32'd0;
     memory[9582] = 32'd0;
     memory[9583] = 32'd0;
     memory[9584] = 32'd0;
     memory[9585] = 32'd1;
     memory[9586] = 32'd0;
     memory[9587] = 32'd1;
     memory[9588] = 32'd1;
     memory[9589] = 32'd1;
     memory[9590] = 32'd1;
     memory[9591] = 32'd0;
     memory[9592] = 32'd1;
     memory[9593] = 32'd1;
     memory[9594] = 32'd0;
     memory[9595] = 32'd1;
     memory[9596] = 32'd0;
     memory[9597] = 32'd1;
     memory[9598] = 32'd1;
     memory[9599] = 32'd0;
     memory[9600] = 32'd0;
     memory[9601] = 32'd1;
     memory[9602] = 32'd1;
     memory[9603] = 32'd1;
     memory[9604] = 32'd1;
     memory[9605] = 32'd1;
     memory[9606] = 32'd0;
     memory[9607] = 32'd0;
     memory[9608] = 32'd0;
     memory[9609] = 32'd0;
     memory[9610] = 32'd0;
     memory[9611] = 32'd1;
     memory[9612] = 32'd1;
     memory[9613] = 32'd0;
     memory[9614] = 32'd1;
     memory[9615] = 32'd0;
     memory[9616] = 32'd1;
     memory[9617] = 32'd1;
     memory[9618] = 32'd1;
     memory[9619] = 32'd0;
     memory[9620] = 32'd0;
     memory[9621] = 32'd0;
     memory[9622] = 32'd1;
     memory[9623] = 32'd1;
     memory[9624] = 32'd0;
     memory[9625] = 32'd1;
     memory[9626] = 32'd0;
     memory[9627] = 32'd1;
     memory[9628] = 32'd1;
     memory[9629] = 32'd1;
     memory[9630] = 32'd1;
     memory[9631] = 32'd0;
     memory[9632] = 32'd1;
     memory[9633] = 32'd0;
     memory[9634] = 32'd1;
     memory[9635] = 32'd0;
     memory[9636] = 32'd0;
     memory[9637] = 32'd0;
     memory[9638] = 32'd1;
     memory[9639] = 32'd0;
     memory[9640] = 32'd1;
     memory[9641] = 32'd1;
     memory[9642] = 32'd1;
     memory[9643] = 32'd0;
     memory[9644] = 32'd0;
     memory[9645] = 32'd0;
     memory[9646] = 32'd1;
     memory[9647] = 32'd1;
     memory[9648] = 32'd1;
     memory[9649] = 32'd1;
     memory[9650] = 32'd1;
     memory[9651] = 32'd0;
     memory[9652] = 32'd1;
     memory[9653] = 32'd0;
     memory[9654] = 32'd1;
     memory[9655] = 32'd1;
     memory[9656] = 32'd0;
     memory[9657] = 32'd1;
     memory[9658] = 32'd0;
     memory[9659] = 32'd0;
     memory[9660] = 32'd1;
     memory[9661] = 32'd0;
     memory[9662] = 32'd0;
     memory[9663] = 32'd0;
     memory[9664] = 32'd1;
     memory[9665] = 32'd0;
     memory[9666] = 32'd0;
     memory[9667] = 32'd1;
     memory[9668] = 32'd1;
     memory[9669] = 32'd0;
     memory[9670] = 32'd1;
     memory[9671] = 32'd0;
     memory[9672] = 32'd1;
     memory[9673] = 32'd0;
     memory[9674] = 32'd0;
     memory[9675] = 32'd1;
     memory[9676] = 32'd0;
     memory[9677] = 32'd1;
     memory[9678] = 32'd0;
     memory[9679] = 32'd1;
     memory[9680] = 32'd1;
     memory[9681] = 32'd1;
     memory[9682] = 32'd1;
     memory[9683] = 32'd1;
     memory[9684] = 32'd0;
     memory[9685] = 32'd1;
     memory[9686] = 32'd1;
     memory[9687] = 32'd0;
     memory[9688] = 32'd1;
     memory[9689] = 32'd1;
     memory[9690] = 32'd1;
     memory[9691] = 32'd0;
     memory[9692] = 32'd0;
     memory[9693] = 32'd0;
     memory[9694] = 32'd1;
     memory[9695] = 32'd0;
     memory[9696] = 32'd0;
     memory[9697] = 32'd1;
     memory[9698] = 32'd0;
     memory[9699] = 32'd0;
     memory[9700] = 32'd0;
     memory[9701] = 32'd1;
     memory[9702] = 32'd1;
     memory[9703] = 32'd1;
     memory[9704] = 32'd0;
     memory[9705] = 32'd1;
     memory[9706] = 32'd0;
     memory[9707] = 32'd0;
     memory[9708] = 32'd1;
     memory[9709] = 32'd1;
     memory[9710] = 32'd0;
     memory[9711] = 32'd1;
     memory[9712] = 32'd0;
     memory[9713] = 32'd0;
     memory[9714] = 32'd1;
     memory[9715] = 32'd0;
     memory[9716] = 32'd1;
     memory[9717] = 32'd0;
     memory[9718] = 32'd1;
     memory[9719] = 32'd0;
     memory[9720] = 32'd1;
     memory[9721] = 32'd1;
     memory[9722] = 32'd0;
     memory[9723] = 32'd0;
     memory[9724] = 32'd0;
     memory[9725] = 32'd1;
     memory[9726] = 32'd1;
     memory[9727] = 32'd1;
     memory[9728] = 32'd1;
     memory[9729] = 32'd1;
     memory[9730] = 32'd1;
     memory[9731] = 32'd1;
     memory[9732] = 32'd0;
     memory[9733] = 32'd1;
     memory[9734] = 32'd0;
     memory[9735] = 32'd1;
     memory[9736] = 32'd0;
     memory[9737] = 32'd1;
     memory[9738] = 32'd1;
     memory[9739] = 32'd1;
     memory[9740] = 32'd1;
     memory[9741] = 32'd0;
     memory[9742] = 32'd1;
     memory[9743] = 32'd1;
     memory[9744] = 32'd0;
     memory[9745] = 32'd1;
     memory[9746] = 32'd1;
     memory[9747] = 32'd0;
     memory[9748] = 32'd1;
     memory[9749] = 32'd0;
     memory[9750] = 32'd0;
     memory[9751] = 32'd0;
     memory[9752] = 32'd0;
     memory[9753] = 32'd1;
     memory[9754] = 32'd0;
     memory[9755] = 32'd0;
     memory[9756] = 32'd1;
     memory[9757] = 32'd1;
     memory[9758] = 32'd1;
     memory[9759] = 32'd0;
     memory[9760] = 32'd1;
     memory[9761] = 32'd1;
     memory[9762] = 32'd1;
     memory[9763] = 32'd1;
     memory[9764] = 32'd1;
     memory[9765] = 32'd0;
     memory[9766] = 32'd1;
     memory[9767] = 32'd1;
     memory[9768] = 32'd1;
     memory[9769] = 32'd0;
     memory[9770] = 32'd0;
     memory[9771] = 32'd0;
     memory[9772] = 32'd0;
     memory[9773] = 32'd0;
     memory[9774] = 32'd1;
     memory[9775] = 32'd1;
     memory[9776] = 32'd1;
     memory[9777] = 32'd1;
     memory[9778] = 32'd0;
     memory[9779] = 32'd1;
     memory[9780] = 32'd1;
     memory[9781] = 32'd1;
     memory[9782] = 32'd0;
     memory[9783] = 32'd1;
     memory[9784] = 32'd0;
     memory[9785] = 32'd0;
     memory[9786] = 32'd1;
     memory[9787] = 32'd0;
     memory[9788] = 32'd0;
     memory[9789] = 32'd1;
     memory[9790] = 32'd0;
     memory[9791] = 32'd0;
     memory[9792] = 32'd0;
     memory[9793] = 32'd1;
     memory[9794] = 32'd1;
     memory[9795] = 32'd0;
     memory[9796] = 32'd1;
     memory[9797] = 32'd1;
     memory[9798] = 32'd0;
     memory[9799] = 32'd1;
     memory[9800] = 32'd0;
     memory[9801] = 32'd1;
     memory[9802] = 32'd1;
     memory[9803] = 32'd0;
     memory[9804] = 32'd0;
     memory[9805] = 32'd0;
     memory[9806] = 32'd1;
     memory[9807] = 32'd1;
     memory[9808] = 32'd0;
     memory[9809] = 32'd1;
     memory[9810] = 32'd0;
     memory[9811] = 32'd0;
     memory[9812] = 32'd1;
     memory[9813] = 32'd1;
     memory[9814] = 32'd1;
     memory[9815] = 32'd1;
     memory[9816] = 32'd0;
     memory[9817] = 32'd0;
     memory[9818] = 32'd0;
     memory[9819] = 32'd0;
     memory[9820] = 32'd1;
     memory[9821] = 32'd0;
     memory[9822] = 32'd1;
     memory[9823] = 32'd1;
     memory[9824] = 32'd0;
     memory[9825] = 32'd1;
     memory[9826] = 32'd0;
     memory[9827] = 32'd1;
     memory[9828] = 32'd1;
     memory[9829] = 32'd0;
     memory[9830] = 32'd0;
     memory[9831] = 32'd1;
     memory[9832] = 32'd1;
     memory[9833] = 32'd1;
     memory[9834] = 32'd0;
     memory[9835] = 32'd0;
     memory[9836] = 32'd0;
     memory[9837] = 32'd0;
     memory[9838] = 32'd0;
     memory[9839] = 32'd1;
     memory[9840] = 32'd1;
     memory[9841] = 32'd1;
     memory[9842] = 32'd1;
     memory[9843] = 32'd1;
     memory[9844] = 32'd0;
     memory[9845] = 32'd0;
     memory[9846] = 32'd0;
     memory[9847] = 32'd1;
     memory[9848] = 32'd1;
     memory[9849] = 32'd0;
     memory[9850] = 32'd1;
     memory[9851] = 32'd0;
     memory[9852] = 32'd1;
     memory[9853] = 32'd1;
     memory[9854] = 32'd1;
     memory[9855] = 32'd1;
     memory[9856] = 32'd1;
     memory[9857] = 32'd0;
     memory[9858] = 32'd1;
     memory[9859] = 32'd0;
     memory[9860] = 32'd0;
     memory[9861] = 32'd1;
     memory[9862] = 32'd0;
     memory[9863] = 32'd0;
     memory[9864] = 32'd0;
     memory[9865] = 32'd1;
     memory[9866] = 32'd0;
     memory[9867] = 32'd0;
     memory[9868] = 32'd1;
     memory[9869] = 32'd0;
     memory[9870] = 32'd1;
     memory[9871] = 32'd0;
     memory[9872] = 32'd1;
     memory[9873] = 32'd0;
     memory[9874] = 32'd0;
     memory[9875] = 32'd0;
     memory[9876] = 32'd0;
     memory[9877] = 32'd1;
     memory[9878] = 32'd1;
     memory[9879] = 32'd0;
     memory[9880] = 32'd1;
     memory[9881] = 32'd0;
     memory[9882] = 32'd1;
     memory[9883] = 32'd0;
     memory[9884] = 32'd1;
     memory[9885] = 32'd1;
     memory[9886] = 32'd0;
     memory[9887] = 32'd0;
     memory[9888] = 32'd0;
     memory[9889] = 32'd1;
     memory[9890] = 32'd1;
     memory[9891] = 32'd1;
     memory[9892] = 32'd0;
     memory[9893] = 32'd0;
     memory[9894] = 32'd1;
     memory[9895] = 32'd0;
     memory[9896] = 32'd0;
     memory[9897] = 32'd0;
     memory[9898] = 32'd1;
     memory[9899] = 32'd0;
     memory[9900] = 32'd0;
     memory[9901] = 32'd0;
     memory[9902] = 32'd1;
     memory[9903] = 32'd1;
     memory[9904] = 32'd1;
     memory[9905] = 32'd0;
     memory[9906] = 32'd0;
     memory[9907] = 32'd1;
     memory[9908] = 32'd1;
     memory[9909] = 32'd0;
     memory[9910] = 32'd1;
     memory[9911] = 32'd1;
     memory[9912] = 32'd0;
     memory[9913] = 32'd0;
     memory[9914] = 32'd1;
     memory[9915] = 32'd0;
     memory[9916] = 32'd0;
     memory[9917] = 32'd0;
     memory[9918] = 32'd1;
     memory[9919] = 32'd0;
     memory[9920] = 32'd0;
     memory[9921] = 32'd1;
     memory[9922] = 32'd1;
     memory[9923] = 32'd1;
     memory[9924] = 32'd0;
     memory[9925] = 32'd1;
     memory[9926] = 32'd1;
     memory[9927] = 32'd1;
     memory[9928] = 32'd0;
     memory[9929] = 32'd1;
     memory[9930] = 32'd0;
     memory[9931] = 32'd1;
     memory[9932] = 32'd0;
     memory[9933] = 32'd1;
     memory[9934] = 32'd1;
     memory[9935] = 32'd1;
     memory[9936] = 32'd0;
     memory[9937] = 32'd1;
     memory[9938] = 32'd1;
     memory[9939] = 32'd0;
     memory[9940] = 32'd0;
     memory[9941] = 32'd1;
     memory[9942] = 32'd1;
     memory[9943] = 32'd0;
     memory[9944] = 32'd1;
     memory[9945] = 32'd0;
     memory[9946] = 32'd1;
     memory[9947] = 32'd1;
     memory[9948] = 32'd1;
     memory[9949] = 32'd0;
     memory[9950] = 32'd0;
     memory[9951] = 32'd1;
     memory[9952] = 32'd0;
     memory[9953] = 32'd0;
     memory[9954] = 32'd0;
     memory[9955] = 32'd1;
     memory[9956] = 32'd0;
     memory[9957] = 32'd0;
     memory[9958] = 32'd1;
     memory[9959] = 32'd0;
     memory[9960] = 32'd0;
     memory[9961] = 32'd1;
     memory[9962] = 32'd0;
     memory[9963] = 32'd0;
     memory[9964] = 32'd0;
     memory[9965] = 32'd1;
     memory[9966] = 32'd0;
     memory[9967] = 32'd1;
     memory[9968] = 32'd1;
     memory[9969] = 32'd0;
     memory[9970] = 32'd0;
     memory[9971] = 32'd1;
     memory[9972] = 32'd1;
     memory[9973] = 32'd1;
     memory[9974] = 32'd0;
     memory[9975] = 32'd1;
     memory[9976] = 32'd1;
     memory[9977] = 32'd1;
     memory[9978] = 32'd1;
     memory[9979] = 32'd1;
     memory[9980] = 32'd1;
     memory[9981] = 32'd1;
     memory[9982] = 32'd0;
     memory[9983] = 32'd0;
     memory[9984] = 32'd0;
     memory[9985] = 32'd0;
     memory[9986] = 32'd1;
     memory[9987] = 32'd0;
     memory[9988] = 32'd1;
     memory[9989] = 32'd0;
     memory[9990] = 32'd1;
     memory[9991] = 32'd1;
     memory[9992] = 32'd0;
     memory[9993] = 32'd1;
     memory[9994] = 32'd1;
     memory[9995] = 32'd1;
     memory[9996] = 32'd0;
     memory[9997] = 32'd0;
     memory[9998] = 32'd0;
     memory[9999] = 32'd1;
     memory[10000] = 32'd0;
     memory[10001] = 32'd0;
     memory[10002] = 32'd1;
     memory[10003] = 32'd1;
     memory[10004] = 32'd0;
     memory[10005] = 32'd0;
     memory[10006] = 32'd1;
     memory[10007] = 32'd1;
     memory[10008] = 32'd1;
     memory[10009] = 32'd1;
     memory[10010] = 32'd1;
     memory[10011] = 32'd1;
     memory[10012] = 32'd0;
     memory[10013] = 32'd1;
     memory[10014] = 32'd1;
     memory[10015] = 32'd1;
     memory[10016] = 32'd0;
     memory[10017] = 32'd0;
     memory[10018] = 32'd1;
     memory[10019] = 32'd1;
     memory[10020] = 32'd0;
     memory[10021] = 32'd1;
     memory[10022] = 32'd0;
     memory[10023] = 32'd0;
     memory[10024] = 32'd0;
     memory[10025] = 32'd0;
     memory[10026] = 32'd0;
     memory[10027] = 32'd1;
     memory[10028] = 32'd1;
     memory[10029] = 32'd0;
     memory[10030] = 32'd1;
     memory[10031] = 32'd0;
     memory[10032] = 32'd0;
     memory[10033] = 32'd1;
     memory[10034] = 32'd0;
     memory[10035] = 32'd0;
     memory[10036] = 32'd0;
     memory[10037] = 32'd1;
     memory[10038] = 32'd1;
     memory[10039] = 32'd1;
     memory[10040] = 32'd0;
     memory[10041] = 32'd1;
     memory[10042] = 32'd0;
     memory[10043] = 32'd0;
     memory[10044] = 32'd0;
     memory[10045] = 32'd0;
     memory[10046] = 32'd0;
     memory[10047] = 32'd1;
     memory[10048] = 32'd1;
     memory[10049] = 32'd1;
     memory[10050] = 32'd0;
     memory[10051] = 32'd0;
     memory[10052] = 32'd1;
     memory[10053] = 32'd1;
     memory[10054] = 32'd1;
     memory[10055] = 32'd0;
     memory[10056] = 32'd1;
     memory[10057] = 32'd0;
     memory[10058] = 32'd1;
     memory[10059] = 32'd0;
     memory[10060] = 32'd1;
     memory[10061] = 32'd1;
     memory[10062] = 32'd1;
     memory[10063] = 32'd0;
     memory[10064] = 32'd0;
     memory[10065] = 32'd0;
     memory[10066] = 32'd0;
     memory[10067] = 32'd0;
     memory[10068] = 32'd0;
     memory[10069] = 32'd1;
     memory[10070] = 32'd0;
     memory[10071] = 32'd0;
     memory[10072] = 32'd1;
     memory[10073] = 32'd0;
     memory[10074] = 32'd1;
     memory[10075] = 32'd0;
     memory[10076] = 32'd0;
     memory[10077] = 32'd1;
     memory[10078] = 32'd1;
     memory[10079] = 32'd1;
     memory[10080] = 32'd1;
     memory[10081] = 32'd0;
     memory[10082] = 32'd0;
     memory[10083] = 32'd0;
     memory[10084] = 32'd1;
     memory[10085] = 32'd0;
     memory[10086] = 32'd1;
     memory[10087] = 32'd0;
     memory[10088] = 32'd0;
     memory[10089] = 32'd1;
     memory[10090] = 32'd0;
     memory[10091] = 32'd1;
     memory[10092] = 32'd0;
     memory[10093] = 32'd0;
     memory[10094] = 32'd0;
     memory[10095] = 32'd1;
     memory[10096] = 32'd1;
     memory[10097] = 32'd0;
     memory[10098] = 32'd1;
     memory[10099] = 32'd1;
     memory[10100] = 32'd1;
     memory[10101] = 32'd0;
     memory[10102] = 32'd1;
     memory[10103] = 32'd0;
     memory[10104] = 32'd1;
     memory[10105] = 32'd1;
     memory[10106] = 32'd1;
     memory[10107] = 32'd0;
     memory[10108] = 32'd0;
     memory[10109] = 32'd1;
     memory[10110] = 32'd0;
     memory[10111] = 32'd0;
     memory[10112] = 32'd1;
     memory[10113] = 32'd1;
     memory[10114] = 32'd0;
     memory[10115] = 32'd1;
     memory[10116] = 32'd1;
     memory[10117] = 32'd1;
     memory[10118] = 32'd0;
     memory[10119] = 32'd1;
     memory[10120] = 32'd0;
     memory[10121] = 32'd1;
     memory[10122] = 32'd0;
     memory[10123] = 32'd1;
     memory[10124] = 32'd0;
     memory[10125] = 32'd0;
     memory[10126] = 32'd1;
     memory[10127] = 32'd1;
     memory[10128] = 32'd0;
     memory[10129] = 32'd1;
     memory[10130] = 32'd0;
     memory[10131] = 32'd1;
     memory[10132] = 32'd1;
     memory[10133] = 32'd0;
     memory[10134] = 32'd1;
     memory[10135] = 32'd0;
     memory[10136] = 32'd0;
     memory[10137] = 32'd1;
     memory[10138] = 32'd0;
     memory[10139] = 32'd1;
     memory[10140] = 32'd1;
     memory[10141] = 32'd0;
     memory[10142] = 32'd1;
     memory[10143] = 32'd0;
     memory[10144] = 32'd1;
     memory[10145] = 32'd1;
     memory[10146] = 32'd1;
     memory[10147] = 32'd1;
     memory[10148] = 32'd1;
     memory[10149] = 32'd0;
     memory[10150] = 32'd1;
     memory[10151] = 32'd1;
     memory[10152] = 32'd1;
     memory[10153] = 32'd0;
     memory[10154] = 32'd1;
     memory[10155] = 32'd0;
     memory[10156] = 32'd1;
     memory[10157] = 32'd0;
     memory[10158] = 32'd1;
     memory[10159] = 32'd0;
     memory[10160] = 32'd1;
     memory[10161] = 32'd1;
     memory[10162] = 32'd1;
     memory[10163] = 32'd0;
     memory[10164] = 32'd0;
     memory[10165] = 32'd0;
     memory[10166] = 32'd1;
     memory[10167] = 32'd1;
     memory[10168] = 32'd0;
     memory[10169] = 32'd1;
     memory[10170] = 32'd1;
     memory[10171] = 32'd1;
     memory[10172] = 32'd0;
     memory[10173] = 32'd0;
     memory[10174] = 32'd1;
     memory[10175] = 32'd1;
     memory[10176] = 32'd0;
     memory[10177] = 32'd1;
     memory[10178] = 32'd0;
     memory[10179] = 32'd1;
     memory[10180] = 32'd1;
     memory[10181] = 32'd1;
     memory[10182] = 32'd0;
     memory[10183] = 32'd1;
     memory[10184] = 32'd0;
     memory[10185] = 32'd0;
     memory[10186] = 32'd1;
     memory[10187] = 32'd0;
     memory[10188] = 32'd0;
     memory[10189] = 32'd1;
     memory[10190] = 32'd0;
     memory[10191] = 32'd0;
     memory[10192] = 32'd1;
     memory[10193] = 32'd0;
     memory[10194] = 32'd0;
     memory[10195] = 32'd1;
     memory[10196] = 32'd0;
     memory[10197] = 32'd1;
     memory[10198] = 32'd0;
     memory[10199] = 32'd0;
     memory[10200] = 32'd0;
     memory[10201] = 32'd0;
     memory[10202] = 32'd0;
     memory[10203] = 32'd0;
     memory[10204] = 32'd1;
     memory[10205] = 32'd0;
     memory[10206] = 32'd0;
     memory[10207] = 32'd0;
     memory[10208] = 32'd0;
     memory[10209] = 32'd0;
     memory[10210] = 32'd0;
     memory[10211] = 32'd0;
     memory[10212] = 32'd1;
     memory[10213] = 32'd1;
     memory[10214] = 32'd1;
     memory[10215] = 32'd1;
     memory[10216] = 32'd1;
     memory[10217] = 32'd1;
     memory[10218] = 32'd1;
     memory[10219] = 32'd1;
     memory[10220] = 32'd1;
     memory[10221] = 32'd1;
     memory[10222] = 32'd0;
     memory[10223] = 32'd1;
     memory[10224] = 32'd1;
     memory[10225] = 32'd1;
     memory[10226] = 32'd1;
     memory[10227] = 32'd0;
     memory[10228] = 32'd1;
     memory[10229] = 32'd0;
     memory[10230] = 32'd0;
     memory[10231] = 32'd1;
     memory[10232] = 32'd0;
     memory[10233] = 32'd0;
     memory[10234] = 32'd0;
     memory[10235] = 32'd0;
     memory[10236] = 32'd0;
     memory[10237] = 32'd0;
     memory[10238] = 32'd1;
     memory[10239] = 32'd0;
     memory[10240] = 32'd0;
     memory[10241] = 32'd0;
     memory[10242] = 32'd0;
     memory[10243] = 32'd0;
     memory[10244] = 32'd1;
     memory[10245] = 32'd0;
     memory[10246] = 32'd1;
     memory[10247] = 32'd0;
     memory[10248] = 32'd0;
     memory[10249] = 32'd0;
     memory[10250] = 32'd0;
     memory[10251] = 32'd0;
     memory[10252] = 32'd0;
     memory[10253] = 32'd0;
     memory[10254] = 32'd1;
     memory[10255] = 32'd1;
     memory[10256] = 32'd1;
     memory[10257] = 32'd0;
     memory[10258] = 32'd1;
     memory[10259] = 32'd0;
     memory[10260] = 32'd1;
     memory[10261] = 32'd1;
     memory[10262] = 32'd1;
     memory[10263] = 32'd1;
     memory[10264] = 32'd1;
     memory[10265] = 32'd1;
     memory[10266] = 32'd1;
     memory[10267] = 32'd0;
     memory[10268] = 32'd1;
     memory[10269] = 32'd1;
     memory[10270] = 32'd0;
     memory[10271] = 32'd1;
     memory[10272] = 32'd1;
     memory[10273] = 32'd0;
     memory[10274] = 32'd0;
     memory[10275] = 32'd1;
     memory[10276] = 32'd0;
     memory[10277] = 32'd1;
     memory[10278] = 32'd0;
     memory[10279] = 32'd1;
     memory[10280] = 32'd0;
     memory[10281] = 32'd1;
     memory[10282] = 32'd0;
     memory[10283] = 32'd1;
     memory[10284] = 32'd0;
     memory[10285] = 32'd0;
     memory[10286] = 32'd1;
     memory[10287] = 32'd1;
     memory[10288] = 32'd0;
     memory[10289] = 32'd1;
     memory[10290] = 32'd1;
     memory[10291] = 32'd0;
     memory[10292] = 32'd1;
     memory[10293] = 32'd1;
     memory[10294] = 32'd1;
     memory[10295] = 32'd1;
     memory[10296] = 32'd1;
     memory[10297] = 32'd1;
     memory[10298] = 32'd1;
     memory[10299] = 32'd0;
     memory[10300] = 32'd1;
     memory[10301] = 32'd0;
     memory[10302] = 32'd1;
     memory[10303] = 32'd1;
     memory[10304] = 32'd0;
     memory[10305] = 32'd0;
     memory[10306] = 32'd1;
     memory[10307] = 32'd0;
     memory[10308] = 32'd1;
     memory[10309] = 32'd1;
     memory[10310] = 32'd1;
     memory[10311] = 32'd0;
     memory[10312] = 32'd1;
     memory[10313] = 32'd0;
     memory[10314] = 32'd1;
     memory[10315] = 32'd0;
     memory[10316] = 32'd1;
     memory[10317] = 32'd0;
     memory[10318] = 32'd1;
     memory[10319] = 32'd1;
     memory[10320] = 32'd0;
     memory[10321] = 32'd0;
     memory[10322] = 32'd1;
     memory[10323] = 32'd1;
     memory[10324] = 32'd1;
     memory[10325] = 32'd0;
     memory[10326] = 32'd1;
     memory[10327] = 32'd1;
     memory[10328] = 32'd0;
     memory[10329] = 32'd0;
     memory[10330] = 32'd1;
     memory[10331] = 32'd1;
     memory[10332] = 32'd1;
     memory[10333] = 32'd1;
     memory[10334] = 32'd0;
     memory[10335] = 32'd0;
     memory[10336] = 32'd0;
     memory[10337] = 32'd0;
     memory[10338] = 32'd0;
     memory[10339] = 32'd0;
     memory[10340] = 32'd0;
     memory[10341] = 32'd1;
     memory[10342] = 32'd0;
     memory[10343] = 32'd1;
     memory[10344] = 32'd1;
     memory[10345] = 32'd0;
     memory[10346] = 32'd0;
     memory[10347] = 32'd0;
     memory[10348] = 32'd1;
     memory[10349] = 32'd0;
     memory[10350] = 32'd0;
     memory[10351] = 32'd1;
     memory[10352] = 32'd0;
     memory[10353] = 32'd1;
     memory[10354] = 32'd1;
     memory[10355] = 32'd0;
     memory[10356] = 32'd0;
     memory[10357] = 32'd1;
     memory[10358] = 32'd0;
     memory[10359] = 32'd0;
     memory[10360] = 32'd0;
     memory[10361] = 32'd1;
     memory[10362] = 32'd0;
     memory[10363] = 32'd1;
     memory[10364] = 32'd1;
     memory[10365] = 32'd1;
     memory[10366] = 32'd1;
     memory[10367] = 32'd0;
     memory[10368] = 32'd0;
     memory[10369] = 32'd1;
     memory[10370] = 32'd1;
     memory[10371] = 32'd0;
     memory[10372] = 32'd1;
     memory[10373] = 32'd1;
     memory[10374] = 32'd1;
     memory[10375] = 32'd0;
     memory[10376] = 32'd0;
     memory[10377] = 32'd0;
     memory[10378] = 32'd1;
     memory[10379] = 32'd0;
     memory[10380] = 32'd0;
     memory[10381] = 32'd0;
     memory[10382] = 32'd0;
     memory[10383] = 32'd1;
     memory[10384] = 32'd1;
     memory[10385] = 32'd1;
     memory[10386] = 32'd1;
     memory[10387] = 32'd0;
     memory[10388] = 32'd0;
     memory[10389] = 32'd0;
     memory[10390] = 32'd0;
     memory[10391] = 32'd0;
     memory[10392] = 32'd1;
     memory[10393] = 32'd1;
     memory[10394] = 32'd0;
     memory[10395] = 32'd0;
     memory[10396] = 32'd1;
     memory[10397] = 32'd1;
     memory[10398] = 32'd1;
     memory[10399] = 32'd0;
     memory[10400] = 32'd0;
     memory[10401] = 32'd0;
     memory[10402] = 32'd1;
     memory[10403] = 32'd1;
     memory[10404] = 32'd1;
     memory[10405] = 32'd1;
     memory[10406] = 32'd0;
     memory[10407] = 32'd0;
     memory[10408] = 32'd1;
     memory[10409] = 32'd0;
     memory[10410] = 32'd0;
     memory[10411] = 32'd0;
     memory[10412] = 32'd1;
     memory[10413] = 32'd1;
     memory[10414] = 32'd1;
     memory[10415] = 32'd0;
     memory[10416] = 32'd0;
     memory[10417] = 32'd0;
     memory[10418] = 32'd1;
     memory[10419] = 32'd1;
     memory[10420] = 32'd0;
     memory[10421] = 32'd1;
     memory[10422] = 32'd1;
     memory[10423] = 32'd1;
     memory[10424] = 32'd0;
     memory[10425] = 32'd1;
     memory[10426] = 32'd0;
     memory[10427] = 32'd1;
     memory[10428] = 32'd1;
     memory[10429] = 32'd1;
     memory[10430] = 32'd1;
     memory[10431] = 32'd0;
     memory[10432] = 32'd0;
     memory[10433] = 32'd0;
     memory[10434] = 32'd1;
     memory[10435] = 32'd1;
     memory[10436] = 32'd0;
     memory[10437] = 32'd1;
     memory[10438] = 32'd0;
     memory[10439] = 32'd1;
     memory[10440] = 32'd0;
     memory[10441] = 32'd1;
     memory[10442] = 32'd1;
     memory[10443] = 32'd1;
     memory[10444] = 32'd0;
     memory[10445] = 32'd1;
     memory[10446] = 32'd0;
     memory[10447] = 32'd0;
     memory[10448] = 32'd1;
     memory[10449] = 32'd0;
     memory[10450] = 32'd1;
     memory[10451] = 32'd1;
     memory[10452] = 32'd1;
     memory[10453] = 32'd1;
     memory[10454] = 32'd0;
     memory[10455] = 32'd0;
     memory[10456] = 32'd0;
     memory[10457] = 32'd1;
     memory[10458] = 32'd1;
     memory[10459] = 32'd1;
     memory[10460] = 32'd0;
     memory[10461] = 32'd0;
     memory[10462] = 32'd1;
     memory[10463] = 32'd0;
     memory[10464] = 32'd0;
     memory[10465] = 32'd1;
     memory[10466] = 32'd0;
     memory[10467] = 32'd1;
     memory[10468] = 32'd0;
     memory[10469] = 32'd0;
     memory[10470] = 32'd1;
     memory[10471] = 32'd0;
     memory[10472] = 32'd1;
     memory[10473] = 32'd1;
     memory[10474] = 32'd0;
     memory[10475] = 32'd0;
     memory[10476] = 32'd0;
     memory[10477] = 32'd0;
     memory[10478] = 32'd1;
     memory[10479] = 32'd0;
     memory[10480] = 32'd1;
     memory[10481] = 32'd0;
     memory[10482] = 32'd0;
     memory[10483] = 32'd0;
     memory[10484] = 32'd0;
     memory[10485] = 32'd1;
     memory[10486] = 32'd1;
     memory[10487] = 32'd1;
     memory[10488] = 32'd0;
     memory[10489] = 32'd0;
     memory[10490] = 32'd1;
     memory[10491] = 32'd1;
     memory[10492] = 32'd0;
     memory[10493] = 32'd0;
     memory[10494] = 32'd0;
     memory[10495] = 32'd1;
     memory[10496] = 32'd1;
     memory[10497] = 32'd0;
     memory[10498] = 32'd1;
     memory[10499] = 32'd1;
     memory[10500] = 32'd0;
     memory[10501] = 32'd1;
     memory[10502] = 32'd0;
     memory[10503] = 32'd0;
     memory[10504] = 32'd1;
     memory[10505] = 32'd0;
     memory[10506] = 32'd0;
     memory[10507] = 32'd0;
     memory[10508] = 32'd0;
     memory[10509] = 32'd1;
     memory[10510] = 32'd1;
     memory[10511] = 32'd0;
     memory[10512] = 32'd0;
     memory[10513] = 32'd1;
     memory[10514] = 32'd0;
     memory[10515] = 32'd0;
     memory[10516] = 32'd1;
     memory[10517] = 32'd0;
     memory[10518] = 32'd0;
     memory[10519] = 32'd0;
     memory[10520] = 32'd1;
     memory[10521] = 32'd0;
     memory[10522] = 32'd0;
     memory[10523] = 32'd1;
     memory[10524] = 32'd0;
     memory[10525] = 32'd1;
     memory[10526] = 32'd0;
     memory[10527] = 32'd0;
     memory[10528] = 32'd0;
     memory[10529] = 32'd1;
     memory[10530] = 32'd1;
     memory[10531] = 32'd0;
     memory[10532] = 32'd0;
     memory[10533] = 32'd1;
     memory[10534] = 32'd1;
     memory[10535] = 32'd1;
     memory[10536] = 32'd1;
     memory[10537] = 32'd0;
     memory[10538] = 32'd1;
     memory[10539] = 32'd1;
     memory[10540] = 32'd0;
     memory[10541] = 32'd0;
     memory[10542] = 32'd1;
     memory[10543] = 32'd0;
     memory[10544] = 32'd1;
     memory[10545] = 32'd1;
     memory[10546] = 32'd0;
     memory[10547] = 32'd0;
     memory[10548] = 32'd0;
     memory[10549] = 32'd1;
     memory[10550] = 32'd0;
     memory[10551] = 32'd1;
     memory[10552] = 32'd0;
     memory[10553] = 32'd1;
     memory[10554] = 32'd0;
     memory[10555] = 32'd0;
     memory[10556] = 32'd0;
     memory[10557] = 32'd1;
     memory[10558] = 32'd1;
     memory[10559] = 32'd0;
     memory[10560] = 32'd0;
     memory[10561] = 32'd1;
     memory[10562] = 32'd1;
     memory[10563] = 32'd0;
     memory[10564] = 32'd1;
     memory[10565] = 32'd0;
     memory[10566] = 32'd0;
     memory[10567] = 32'd0;
     memory[10568] = 32'd0;
     memory[10569] = 32'd0;
     memory[10570] = 32'd1;
     memory[10571] = 32'd0;
     memory[10572] = 32'd1;
     memory[10573] = 32'd0;
     memory[10574] = 32'd0;
     memory[10575] = 32'd1;
     memory[10576] = 32'd0;
     memory[10577] = 32'd0;
     memory[10578] = 32'd1;
     memory[10579] = 32'd0;
     memory[10580] = 32'd0;
     memory[10581] = 32'd1;
     memory[10582] = 32'd0;
     memory[10583] = 32'd1;
     memory[10584] = 32'd1;
     memory[10585] = 32'd1;
     memory[10586] = 32'd1;
     memory[10587] = 32'd1;
     memory[10588] = 32'd1;
     memory[10589] = 32'd1;
     memory[10590] = 32'd1;
     memory[10591] = 32'd1;
     memory[10592] = 32'd1;
     memory[10593] = 32'd1;
     memory[10594] = 32'd1;
     memory[10595] = 32'd0;
     memory[10596] = 32'd1;
     memory[10597] = 32'd1;
     memory[10598] = 32'd1;
     memory[10599] = 32'd1;
     memory[10600] = 32'd0;
     memory[10601] = 32'd0;
     memory[10602] = 32'd0;
     memory[10603] = 32'd0;
     memory[10604] = 32'd1;
     memory[10605] = 32'd1;
     memory[10606] = 32'd1;
     memory[10607] = 32'd0;
     memory[10608] = 32'd1;
     memory[10609] = 32'd0;
     memory[10610] = 32'd0;
     memory[10611] = 32'd1;
     memory[10612] = 32'd1;
     memory[10613] = 32'd0;
     memory[10614] = 32'd1;
     memory[10615] = 32'd1;
     memory[10616] = 32'd1;
     memory[10617] = 32'd0;
     memory[10618] = 32'd0;
     memory[10619] = 32'd0;
     memory[10620] = 32'd0;
     memory[10621] = 32'd0;
     memory[10622] = 32'd0;
     memory[10623] = 32'd0;
     memory[10624] = 32'd1;
     memory[10625] = 32'd1;
     memory[10626] = 32'd1;
     memory[10627] = 32'd1;
     memory[10628] = 32'd0;
     memory[10629] = 32'd1;
     memory[10630] = 32'd0;
     memory[10631] = 32'd0;
     memory[10632] = 32'd0;
     memory[10633] = 32'd0;
     memory[10634] = 32'd0;
     memory[10635] = 32'd1;
     memory[10636] = 32'd1;
     memory[10637] = 32'd0;
     memory[10638] = 32'd0;
     memory[10639] = 32'd0;
     memory[10640] = 32'd0;
     memory[10641] = 32'd0;
     memory[10642] = 32'd1;
     memory[10643] = 32'd1;
     memory[10644] = 32'd0;
     memory[10645] = 32'd1;
     memory[10646] = 32'd0;
     memory[10647] = 32'd0;
     memory[10648] = 32'd1;
     memory[10649] = 32'd1;
     memory[10650] = 32'd0;
     memory[10651] = 32'd1;
     memory[10652] = 32'd1;
     memory[10653] = 32'd0;
     memory[10654] = 32'd1;
     memory[10655] = 32'd0;
     memory[10656] = 32'd1;
     memory[10657] = 32'd1;
     memory[10658] = 32'd0;
     memory[10659] = 32'd1;
     memory[10660] = 32'd0;
     memory[10661] = 32'd0;
     memory[10662] = 32'd1;
     memory[10663] = 32'd1;
     memory[10664] = 32'd1;
     memory[10665] = 32'd1;
     memory[10666] = 32'd1;
     memory[10667] = 32'd1;
     memory[10668] = 32'd0;
     memory[10669] = 32'd1;
     memory[10670] = 32'd1;
     memory[10671] = 32'd1;
     memory[10672] = 32'd0;
     memory[10673] = 32'd0;
     memory[10674] = 32'd1;
     memory[10675] = 32'd1;
     memory[10676] = 32'd1;
     memory[10677] = 32'd0;
     memory[10678] = 32'd1;
     memory[10679] = 32'd1;
     memory[10680] = 32'd1;
     memory[10681] = 32'd0;
     memory[10682] = 32'd0;
     memory[10683] = 32'd0;
     memory[10684] = 32'd0;
     memory[10685] = 32'd0;
     memory[10686] = 32'd0;
     memory[10687] = 32'd0;
     memory[10688] = 32'd1;
     memory[10689] = 32'd1;
     memory[10690] = 32'd1;
     memory[10691] = 32'd1;
     memory[10692] = 32'd1;
     memory[10693] = 32'd0;
     memory[10694] = 32'd0;
     memory[10695] = 32'd0;
     memory[10696] = 32'd0;
     memory[10697] = 32'd1;
     memory[10698] = 32'd1;
     memory[10699] = 32'd0;
     memory[10700] = 32'd0;
     memory[10701] = 32'd1;
     memory[10702] = 32'd0;
     memory[10703] = 32'd1;
     memory[10704] = 32'd1;
     memory[10705] = 32'd1;
     memory[10706] = 32'd1;
     memory[10707] = 32'd0;
     memory[10708] = 32'd1;
     memory[10709] = 32'd1;
     memory[10710] = 32'd0;
     memory[10711] = 32'd0;
     memory[10712] = 32'd1;
     memory[10713] = 32'd0;
     memory[10714] = 32'd0;
     memory[10715] = 32'd1;
     memory[10716] = 32'd0;
     memory[10717] = 32'd1;
     memory[10718] = 32'd1;
     memory[10719] = 32'd1;
     memory[10720] = 32'd1;
     memory[10721] = 32'd0;
     memory[10722] = 32'd1;
     memory[10723] = 32'd0;
     memory[10724] = 32'd1;
     memory[10725] = 32'd0;
     memory[10726] = 32'd0;
     memory[10727] = 32'd1;
     memory[10728] = 32'd1;
     memory[10729] = 32'd0;
     memory[10730] = 32'd0;
     memory[10731] = 32'd0;
     memory[10732] = 32'd1;
     memory[10733] = 32'd0;
     memory[10734] = 32'd1;
     memory[10735] = 32'd1;
     memory[10736] = 32'd1;
     memory[10737] = 32'd0;
     memory[10738] = 32'd1;
     memory[10739] = 32'd0;
     memory[10740] = 32'd1;
     memory[10741] = 32'd1;
     memory[10742] = 32'd0;
     memory[10743] = 32'd0;
     memory[10744] = 32'd0;
     memory[10745] = 32'd0;
     memory[10746] = 32'd0;
     memory[10747] = 32'd0;
     memory[10748] = 32'd1;
     memory[10749] = 32'd1;
     memory[10750] = 32'd0;
     memory[10751] = 32'd1;
     memory[10752] = 32'd1;
     memory[10753] = 32'd0;
     memory[10754] = 32'd0;
     memory[10755] = 32'd1;
     memory[10756] = 32'd1;
     memory[10757] = 32'd0;
     memory[10758] = 32'd0;
     memory[10759] = 32'd1;
     memory[10760] = 32'd1;
     memory[10761] = 32'd0;
     memory[10762] = 32'd1;
     memory[10763] = 32'd1;
     memory[10764] = 32'd1;
     memory[10765] = 32'd1;
     memory[10766] = 32'd0;
     memory[10767] = 32'd1;
     memory[10768] = 32'd0;
     memory[10769] = 32'd1;
     memory[10770] = 32'd0;
     memory[10771] = 32'd0;
     memory[10772] = 32'd1;
     memory[10773] = 32'd0;
     memory[10774] = 32'd1;
     memory[10775] = 32'd1;
     memory[10776] = 32'd1;
     memory[10777] = 32'd1;
     memory[10778] = 32'd0;
     memory[10779] = 32'd1;
     memory[10780] = 32'd0;
     memory[10781] = 32'd0;
     memory[10782] = 32'd0;
     memory[10783] = 32'd1;
     memory[10784] = 32'd0;
     memory[10785] = 32'd1;
     memory[10786] = 32'd0;
     memory[10787] = 32'd1;
     memory[10788] = 32'd0;
     memory[10789] = 32'd1;
     memory[10790] = 32'd0;
     memory[10791] = 32'd0;
     memory[10792] = 32'd0;
     memory[10793] = 32'd0;
     memory[10794] = 32'd0;
     memory[10795] = 32'd1;
     memory[10796] = 32'd1;
     memory[10797] = 32'd1;
     memory[10798] = 32'd1;
     memory[10799] = 32'd1;
     memory[10800] = 32'd1;
     memory[10801] = 32'd1;
     memory[10802] = 32'd0;
     memory[10803] = 32'd0;
     memory[10804] = 32'd1;
     memory[10805] = 32'd0;
     memory[10806] = 32'd0;
     memory[10807] = 32'd0;
     memory[10808] = 32'd1;
     memory[10809] = 32'd0;
     memory[10810] = 32'd0;
     memory[10811] = 32'd0;
     memory[10812] = 32'd0;
     memory[10813] = 32'd1;
     memory[10814] = 32'd1;
     memory[10815] = 32'd0;
     memory[10816] = 32'd1;
     memory[10817] = 32'd0;
     memory[10818] = 32'd0;
     memory[10819] = 32'd1;
     memory[10820] = 32'd1;
     memory[10821] = 32'd1;
     memory[10822] = 32'd0;
     memory[10823] = 32'd1;
     memory[10824] = 32'd0;
     memory[10825] = 32'd1;
     memory[10826] = 32'd1;
     memory[10827] = 32'd0;
     memory[10828] = 32'd1;
     memory[10829] = 32'd0;
     memory[10830] = 32'd0;
     memory[10831] = 32'd1;
     memory[10832] = 32'd1;
     memory[10833] = 32'd0;
     memory[10834] = 32'd0;
     memory[10835] = 32'd1;
     memory[10836] = 32'd1;
     memory[10837] = 32'd1;
     memory[10838] = 32'd0;
     memory[10839] = 32'd1;
     memory[10840] = 32'd1;
     memory[10841] = 32'd1;
     memory[10842] = 32'd0;
     memory[10843] = 32'd1;
     memory[10844] = 32'd1;
     memory[10845] = 32'd1;
     memory[10846] = 32'd1;
     memory[10847] = 32'd0;
     memory[10848] = 32'd0;
     memory[10849] = 32'd0;
     memory[10850] = 32'd0;
     memory[10851] = 32'd1;
     memory[10852] = 32'd1;
     memory[10853] = 32'd1;
     memory[10854] = 32'd0;
     memory[10855] = 32'd0;
     memory[10856] = 32'd1;
     memory[10857] = 32'd1;
     memory[10858] = 32'd1;
     memory[10859] = 32'd1;
     memory[10860] = 32'd0;
     memory[10861] = 32'd0;
     memory[10862] = 32'd1;
     memory[10863] = 32'd0;
     memory[10864] = 32'd0;
     memory[10865] = 32'd0;
     memory[10866] = 32'd1;
     memory[10867] = 32'd1;
     memory[10868] = 32'd1;
     memory[10869] = 32'd1;
     memory[10870] = 32'd1;
     memory[10871] = 32'd1;
     memory[10872] = 32'd1;
     memory[10873] = 32'd1;
     memory[10874] = 32'd0;
     memory[10875] = 32'd0;
     memory[10876] = 32'd0;
     memory[10877] = 32'd1;
     memory[10878] = 32'd0;
     memory[10879] = 32'd0;
     memory[10880] = 32'd1;
     memory[10881] = 32'd0;
     memory[10882] = 32'd1;
     memory[10883] = 32'd0;
     memory[10884] = 32'd0;
     memory[10885] = 32'd1;
     memory[10886] = 32'd0;
     memory[10887] = 32'd1;
     memory[10888] = 32'd1;
     memory[10889] = 32'd0;
     memory[10890] = 32'd0;
     memory[10891] = 32'd0;
     memory[10892] = 32'd0;
     memory[10893] = 32'd0;
     memory[10894] = 32'd1;
     memory[10895] = 32'd1;
     memory[10896] = 32'd1;
     memory[10897] = 32'd1;
     memory[10898] = 32'd0;
     memory[10899] = 32'd0;
     memory[10900] = 32'd0;
     memory[10901] = 32'd0;
     memory[10902] = 32'd1;
     memory[10903] = 32'd1;
     memory[10904] = 32'd0;
     memory[10905] = 32'd0;
     memory[10906] = 32'd1;
     memory[10907] = 32'd1;
     memory[10908] = 32'd1;
     memory[10909] = 32'd1;
     memory[10910] = 32'd0;
     memory[10911] = 32'd1;
     memory[10912] = 32'd1;
     memory[10913] = 32'd1;
     memory[10914] = 32'd0;
     memory[10915] = 32'd1;
     memory[10916] = 32'd0;
     memory[10917] = 32'd0;
     memory[10918] = 32'd0;
     memory[10919] = 32'd0;
     memory[10920] = 32'd0;
     memory[10921] = 32'd0;
     memory[10922] = 32'd1;
     memory[10923] = 32'd0;
     memory[10924] = 32'd0;
     memory[10925] = 32'd1;
     memory[10926] = 32'd1;
     memory[10927] = 32'd0;
     memory[10928] = 32'd0;
     memory[10929] = 32'd1;
     memory[10930] = 32'd1;
     memory[10931] = 32'd0;
     memory[10932] = 32'd0;
     memory[10933] = 32'd0;
     memory[10934] = 32'd1;
     memory[10935] = 32'd1;
     memory[10936] = 32'd0;
     memory[10937] = 32'd1;
     memory[10938] = 32'd1;
     memory[10939] = 32'd0;
     memory[10940] = 32'd1;
     memory[10941] = 32'd1;
     memory[10942] = 32'd1;
     memory[10943] = 32'd1;
     memory[10944] = 32'd1;
     memory[10945] = 32'd0;
     memory[10946] = 32'd1;
     memory[10947] = 32'd1;
     memory[10948] = 32'd1;
     memory[10949] = 32'd0;
     memory[10950] = 32'd1;
     memory[10951] = 32'd1;
     memory[10952] = 32'd0;
     memory[10953] = 32'd0;
     memory[10954] = 32'd0;
     memory[10955] = 32'd1;
     memory[10956] = 32'd1;
     memory[10957] = 32'd1;
     memory[10958] = 32'd0;
     memory[10959] = 32'd0;
     memory[10960] = 32'd0;
     memory[10961] = 32'd1;
     memory[10962] = 32'd1;
     memory[10963] = 32'd0;
     memory[10964] = 32'd0;
     memory[10965] = 32'd1;
     memory[10966] = 32'd0;
     memory[10967] = 32'd1;
     memory[10968] = 32'd1;
     memory[10969] = 32'd1;
     memory[10970] = 32'd1;
     memory[10971] = 32'd1;
     memory[10972] = 32'd1;
     memory[10973] = 32'd1;
     memory[10974] = 32'd1;
     memory[10975] = 32'd1;
     memory[10976] = 32'd0;
     memory[10977] = 32'd0;
     memory[10978] = 32'd1;
     memory[10979] = 32'd1;
     memory[10980] = 32'd1;
     memory[10981] = 32'd1;
     memory[10982] = 32'd1;
     memory[10983] = 32'd1;
     memory[10984] = 32'd1;
     memory[10985] = 32'd1;
     memory[10986] = 32'd1;
     memory[10987] = 32'd1;
     memory[10988] = 32'd1;
     memory[10989] = 32'd1;
     memory[10990] = 32'd1;
     memory[10991] = 32'd1;
     memory[10992] = 32'd1;
     memory[10993] = 32'd0;
     memory[10994] = 32'd0;
     memory[10995] = 32'd1;
     memory[10996] = 32'd1;
     memory[10997] = 32'd0;
     memory[10998] = 32'd1;
     memory[10999] = 32'd0;
     memory[11000] = 32'd1;
     memory[11001] = 32'd0;
     memory[11002] = 32'd1;
     memory[11003] = 32'd0;
     memory[11004] = 32'd1;
     memory[11005] = 32'd0;
     memory[11006] = 32'd1;
     memory[11007] = 32'd1;
     memory[11008] = 32'd0;
     memory[11009] = 32'd0;
     memory[11010] = 32'd0;
     memory[11011] = 32'd1;
     memory[11012] = 32'd1;
     memory[11013] = 32'd0;
     memory[11014] = 32'd1;
     memory[11015] = 32'd1;
     memory[11016] = 32'd0;
     memory[11017] = 32'd1;
     memory[11018] = 32'd1;
     memory[11019] = 32'd1;
     memory[11020] = 32'd1;
     memory[11021] = 32'd1;
     memory[11022] = 32'd0;
     memory[11023] = 32'd1;
     memory[11024] = 32'd0;
     memory[11025] = 32'd0;
     memory[11026] = 32'd1;
     memory[11027] = 32'd1;
     memory[11028] = 32'd0;
     memory[11029] = 32'd0;
     memory[11030] = 32'd0;
     memory[11031] = 32'd0;
     memory[11032] = 32'd0;
     memory[11033] = 32'd1;
     memory[11034] = 32'd0;
     memory[11035] = 32'd1;
     memory[11036] = 32'd0;
     memory[11037] = 32'd0;
     memory[11038] = 32'd1;
     memory[11039] = 32'd0;
     memory[11040] = 32'd1;
     memory[11041] = 32'd1;
     memory[11042] = 32'd1;
     memory[11043] = 32'd0;
     memory[11044] = 32'd0;
     memory[11045] = 32'd1;
     memory[11046] = 32'd1;
     memory[11047] = 32'd0;
     memory[11048] = 32'd1;
     memory[11049] = 32'd1;
     memory[11050] = 32'd1;
     memory[11051] = 32'd0;
     memory[11052] = 32'd0;
     memory[11053] = 32'd1;
     memory[11054] = 32'd0;
     memory[11055] = 32'd0;
     memory[11056] = 32'd1;
     memory[11057] = 32'd1;
     memory[11058] = 32'd1;
     memory[11059] = 32'd0;
     memory[11060] = 32'd1;
     memory[11061] = 32'd1;
     memory[11062] = 32'd0;
     memory[11063] = 32'd0;
     memory[11064] = 32'd1;
     memory[11065] = 32'd1;
     memory[11066] = 32'd1;
     memory[11067] = 32'd1;
     memory[11068] = 32'd0;
     memory[11069] = 32'd0;
     memory[11070] = 32'd1;
     memory[11071] = 32'd1;
     memory[11072] = 32'd1;
     memory[11073] = 32'd1;
     memory[11074] = 32'd1;
     memory[11075] = 32'd0;
     memory[11076] = 32'd1;
     memory[11077] = 32'd1;
     memory[11078] = 32'd1;
     memory[11079] = 32'd1;
     memory[11080] = 32'd0;
     memory[11081] = 32'd0;
     memory[11082] = 32'd0;
     memory[11083] = 32'd0;
     memory[11084] = 32'd0;
     memory[11085] = 32'd0;
     memory[11086] = 32'd0;
     memory[11087] = 32'd0;
     memory[11088] = 32'd1;
     memory[11089] = 32'd0;
     memory[11090] = 32'd1;
     memory[11091] = 32'd0;
     memory[11092] = 32'd0;
     memory[11093] = 32'd0;
     memory[11094] = 32'd1;
     memory[11095] = 32'd1;
     memory[11096] = 32'd0;
     memory[11097] = 32'd1;
     memory[11098] = 32'd1;
     memory[11099] = 32'd0;
     memory[11100] = 32'd1;
     memory[11101] = 32'd1;
     memory[11102] = 32'd1;
     memory[11103] = 32'd0;
     memory[11104] = 32'd0;
     memory[11105] = 32'd1;
     memory[11106] = 32'd0;
     memory[11107] = 32'd0;
     memory[11108] = 32'd1;
     memory[11109] = 32'd1;
     memory[11110] = 32'd1;
     memory[11111] = 32'd0;
     memory[11112] = 32'd0;
     memory[11113] = 32'd0;
     memory[11114] = 32'd1;
     memory[11115] = 32'd0;
     memory[11116] = 32'd1;
     memory[11117] = 32'd1;
     memory[11118] = 32'd0;
     memory[11119] = 32'd1;
     memory[11120] = 32'd1;
     memory[11121] = 32'd0;
     memory[11122] = 32'd0;
     memory[11123] = 32'd0;
     memory[11124] = 32'd1;
     memory[11125] = 32'd1;
     memory[11126] = 32'd1;
     memory[11127] = 32'd0;
     memory[11128] = 32'd0;
     memory[11129] = 32'd1;
     memory[11130] = 32'd1;
     memory[11131] = 32'd0;
     memory[11132] = 32'd1;
     memory[11133] = 32'd1;
     memory[11134] = 32'd0;
     memory[11135] = 32'd1;
     memory[11136] = 32'd1;
     memory[11137] = 32'd1;
     memory[11138] = 32'd0;
     memory[11139] = 32'd1;
     memory[11140] = 32'd1;
     memory[11141] = 32'd0;
     memory[11142] = 32'd1;
     memory[11143] = 32'd1;
     memory[11144] = 32'd1;
     memory[11145] = 32'd0;
     memory[11146] = 32'd0;
     memory[11147] = 32'd1;
     memory[11148] = 32'd1;
     memory[11149] = 32'd0;
     memory[11150] = 32'd1;
     memory[11151] = 32'd1;
     memory[11152] = 32'd0;
     memory[11153] = 32'd0;
     memory[11154] = 32'd0;
     memory[11155] = 32'd0;
     memory[11156] = 32'd1;
     memory[11157] = 32'd0;
     memory[11158] = 32'd0;
     memory[11159] = 32'd1;
     memory[11160] = 32'd0;
     memory[11161] = 32'd1;
     memory[11162] = 32'd0;
     memory[11163] = 32'd0;
     memory[11164] = 32'd1;
     memory[11165] = 32'd0;
     memory[11166] = 32'd1;
     memory[11167] = 32'd1;
     memory[11168] = 32'd1;
     memory[11169] = 32'd1;
     memory[11170] = 32'd0;
     memory[11171] = 32'd0;
     memory[11172] = 32'd0;
     memory[11173] = 32'd0;
     memory[11174] = 32'd0;
     memory[11175] = 32'd1;
     memory[11176] = 32'd0;
     memory[11177] = 32'd1;
     memory[11178] = 32'd0;
     memory[11179] = 32'd1;
     memory[11180] = 32'd0;
     memory[11181] = 32'd1;
     memory[11182] = 32'd1;
     memory[11183] = 32'd0;
     memory[11184] = 32'd0;
     memory[11185] = 32'd1;
     memory[11186] = 32'd1;
     memory[11187] = 32'd0;
     memory[11188] = 32'd1;
     memory[11189] = 32'd1;
     memory[11190] = 32'd1;
     memory[11191] = 32'd0;
     memory[11192] = 32'd1;
     memory[11193] = 32'd1;
     memory[11194] = 32'd0;
     memory[11195] = 32'd1;
     memory[11196] = 32'd1;
     memory[11197] = 32'd1;
     memory[11198] = 32'd0;
     memory[11199] = 32'd0;
     memory[11200] = 32'd0;
     memory[11201] = 32'd1;
     memory[11202] = 32'd1;
     memory[11203] = 32'd1;
     memory[11204] = 32'd0;
     memory[11205] = 32'd0;
     memory[11206] = 32'd0;
     memory[11207] = 32'd0;
     memory[11208] = 32'd1;
     memory[11209] = 32'd1;
     memory[11210] = 32'd1;
     memory[11211] = 32'd1;
     memory[11212] = 32'd1;
     memory[11213] = 32'd1;
     memory[11214] = 32'd1;
     memory[11215] = 32'd0;
     memory[11216] = 32'd1;
     memory[11217] = 32'd1;
     memory[11218] = 32'd0;
     memory[11219] = 32'd1;
     memory[11220] = 32'd0;
     memory[11221] = 32'd0;
     memory[11222] = 32'd0;
     memory[11223] = 32'd0;
     memory[11224] = 32'd1;
     memory[11225] = 32'd0;
     memory[11226] = 32'd1;
     memory[11227] = 32'd0;
     memory[11228] = 32'd0;
     memory[11229] = 32'd1;
     memory[11230] = 32'd0;
     memory[11231] = 32'd1;
     memory[11232] = 32'd0;
     memory[11233] = 32'd0;
     memory[11234] = 32'd0;
     memory[11235] = 32'd1;
     memory[11236] = 32'd1;
     memory[11237] = 32'd1;
     memory[11238] = 32'd0;
     memory[11239] = 32'd1;
     memory[11240] = 32'd0;
     memory[11241] = 32'd0;
     memory[11242] = 32'd1;
     memory[11243] = 32'd1;
     memory[11244] = 32'd1;
     memory[11245] = 32'd1;
     memory[11246] = 32'd1;
     memory[11247] = 32'd0;
     memory[11248] = 32'd0;
     memory[11249] = 32'd1;
     memory[11250] = 32'd1;
     memory[11251] = 32'd0;
     memory[11252] = 32'd1;
     memory[11253] = 32'd0;
     memory[11254] = 32'd1;
     memory[11255] = 32'd0;
     memory[11256] = 32'd1;
     memory[11257] = 32'd0;
     memory[11258] = 32'd1;
     memory[11259] = 32'd1;
     memory[11260] = 32'd0;
     memory[11261] = 32'd1;
     memory[11262] = 32'd0;
     memory[11263] = 32'd0;
     memory[11264] = 32'd1;
     memory[11265] = 32'd1;
     memory[11266] = 32'd1;
     memory[11267] = 32'd0;
     memory[11268] = 32'd1;
     memory[11269] = 32'd1;
     memory[11270] = 32'd1;
     memory[11271] = 32'd0;
     memory[11272] = 32'd0;
     memory[11273] = 32'd1;
     memory[11274] = 32'd0;
     memory[11275] = 32'd1;
     memory[11276] = 32'd1;
     memory[11277] = 32'd0;
     memory[11278] = 32'd0;
     memory[11279] = 32'd0;
     memory[11280] = 32'd1;
     memory[11281] = 32'd0;
     memory[11282] = 32'd0;
     memory[11283] = 32'd1;
     memory[11284] = 32'd1;
     memory[11285] = 32'd0;
     memory[11286] = 32'd0;
     memory[11287] = 32'd1;
     memory[11288] = 32'd1;
     memory[11289] = 32'd1;
     memory[11290] = 32'd1;
     memory[11291] = 32'd0;
     memory[11292] = 32'd0;
     memory[11293] = 32'd0;
     memory[11294] = 32'd1;
     memory[11295] = 32'd1;
     memory[11296] = 32'd1;
     memory[11297] = 32'd0;
     memory[11298] = 32'd0;
     memory[11299] = 32'd1;
     memory[11300] = 32'd0;
     memory[11301] = 32'd0;
     memory[11302] = 32'd0;
     memory[11303] = 32'd1;
     memory[11304] = 32'd1;
     memory[11305] = 32'd0;
     memory[11306] = 32'd0;
     memory[11307] = 32'd1;
     memory[11308] = 32'd1;
     memory[11309] = 32'd1;
     memory[11310] = 32'd1;
     memory[11311] = 32'd1;
     memory[11312] = 32'd1;
     memory[11313] = 32'd1;
     memory[11314] = 32'd0;
     memory[11315] = 32'd1;
     memory[11316] = 32'd1;
     memory[11317] = 32'd0;
     memory[11318] = 32'd1;
     memory[11319] = 32'd1;
     memory[11320] = 32'd0;
     memory[11321] = 32'd0;
     memory[11322] = 32'd0;
     memory[11323] = 32'd0;
     memory[11324] = 32'd0;
     memory[11325] = 32'd1;
     memory[11326] = 32'd0;
     memory[11327] = 32'd1;
     memory[11328] = 32'd1;
     memory[11329] = 32'd1;
     memory[11330] = 32'd1;
     memory[11331] = 32'd0;
     memory[11332] = 32'd0;
     memory[11333] = 32'd0;
     memory[11334] = 32'd0;
     memory[11335] = 32'd0;
     memory[11336] = 32'd1;
     memory[11337] = 32'd1;
     memory[11338] = 32'd1;
     memory[11339] = 32'd1;
     memory[11340] = 32'd0;
     memory[11341] = 32'd1;
     memory[11342] = 32'd1;
     memory[11343] = 32'd0;
     memory[11344] = 32'd1;
     memory[11345] = 32'd1;
     memory[11346] = 32'd0;
     memory[11347] = 32'd0;
     memory[11348] = 32'd1;
     memory[11349] = 32'd1;
     memory[11350] = 32'd0;
     memory[11351] = 32'd1;
     memory[11352] = 32'd1;
     memory[11353] = 32'd1;
     memory[11354] = 32'd0;
     memory[11355] = 32'd1;
     memory[11356] = 32'd1;
     memory[11357] = 32'd0;
     memory[11358] = 32'd1;
     memory[11359] = 32'd1;
     memory[11360] = 32'd1;
     memory[11361] = 32'd1;
     memory[11362] = 32'd0;
     memory[11363] = 32'd1;
     memory[11364] = 32'd1;
     memory[11365] = 32'd0;
     memory[11366] = 32'd1;
     memory[11367] = 32'd0;
     memory[11368] = 32'd1;
     memory[11369] = 32'd1;
     memory[11370] = 32'd0;
     memory[11371] = 32'd1;
     memory[11372] = 32'd1;
     memory[11373] = 32'd0;
     memory[11374] = 32'd1;
     memory[11375] = 32'd0;
     memory[11376] = 32'd1;
     memory[11377] = 32'd1;
     memory[11378] = 32'd0;
     memory[11379] = 32'd1;
     memory[11380] = 32'd1;
     memory[11381] = 32'd1;
     memory[11382] = 32'd0;
     memory[11383] = 32'd1;
     memory[11384] = 32'd1;
     memory[11385] = 32'd1;
     memory[11386] = 32'd0;
     memory[11387] = 32'd0;
     memory[11388] = 32'd1;
     memory[11389] = 32'd1;
     memory[11390] = 32'd0;
     memory[11391] = 32'd1;
     memory[11392] = 32'd0;
     memory[11393] = 32'd0;
     memory[11394] = 32'd1;
     memory[11395] = 32'd0;
     memory[11396] = 32'd1;
     memory[11397] = 32'd0;
     memory[11398] = 32'd0;
     memory[11399] = 32'd0;
     memory[11400] = 32'd1;
     memory[11401] = 32'd1;
     memory[11402] = 32'd0;
     memory[11403] = 32'd1;
     memory[11404] = 32'd0;
     memory[11405] = 32'd1;
     memory[11406] = 32'd0;
     memory[11407] = 32'd1;
     memory[11408] = 32'd1;
     memory[11409] = 32'd0;
     memory[11410] = 32'd1;
     memory[11411] = 32'd1;
     memory[11412] = 32'd1;
     memory[11413] = 32'd1;
     memory[11414] = 32'd1;
     memory[11415] = 32'd0;
     memory[11416] = 32'd0;
     memory[11417] = 32'd1;
     memory[11418] = 32'd1;
     memory[11419] = 32'd0;
     memory[11420] = 32'd0;
     memory[11421] = 32'd0;
     memory[11422] = 32'd0;
     memory[11423] = 32'd1;
     memory[11424] = 32'd0;
     memory[11425] = 32'd1;
     memory[11426] = 32'd1;
     memory[11427] = 32'd0;
     memory[11428] = 32'd0;
     memory[11429] = 32'd1;
     memory[11430] = 32'd0;
     memory[11431] = 32'd1;
     memory[11432] = 32'd0;
     memory[11433] = 32'd0;
     memory[11434] = 32'd1;
     memory[11435] = 32'd0;
     memory[11436] = 32'd0;
     memory[11437] = 32'd0;
     memory[11438] = 32'd1;
     memory[11439] = 32'd1;
     memory[11440] = 32'd0;
     memory[11441] = 32'd0;
     memory[11442] = 32'd0;
     memory[11443] = 32'd0;
     memory[11444] = 32'd0;
     memory[11445] = 32'd0;
     memory[11446] = 32'd1;
     memory[11447] = 32'd0;
     memory[11448] = 32'd0;
     memory[11449] = 32'd0;
     memory[11450] = 32'd1;
     memory[11451] = 32'd1;
     memory[11452] = 32'd0;
     memory[11453] = 32'd1;
     memory[11454] = 32'd1;
     memory[11455] = 32'd0;
     memory[11456] = 32'd0;
     memory[11457] = 32'd1;
     memory[11458] = 32'd0;
     memory[11459] = 32'd0;
     memory[11460] = 32'd0;
     memory[11461] = 32'd1;
     memory[11462] = 32'd0;
     memory[11463] = 32'd0;
     memory[11464] = 32'd0;
     memory[11465] = 32'd0;
     memory[11466] = 32'd0;
     memory[11467] = 32'd1;
     memory[11468] = 32'd0;
     memory[11469] = 32'd1;
     memory[11470] = 32'd1;
     memory[11471] = 32'd1;
     memory[11472] = 32'd0;
     memory[11473] = 32'd1;
     memory[11474] = 32'd0;
     memory[11475] = 32'd0;
     memory[11476] = 32'd1;
     memory[11477] = 32'd1;
     memory[11478] = 32'd0;
     memory[11479] = 32'd0;
     memory[11480] = 32'd0;
     memory[11481] = 32'd1;
     memory[11482] = 32'd1;
     memory[11483] = 32'd1;
     memory[11484] = 32'd0;
     memory[11485] = 32'd1;
     memory[11486] = 32'd0;
     memory[11487] = 32'd0;
     memory[11488] = 32'd0;
     memory[11489] = 32'd0;
     memory[11490] = 32'd0;
     memory[11491] = 32'd0;
     memory[11492] = 32'd0;
     memory[11493] = 32'd1;
     memory[11494] = 32'd0;
     memory[11495] = 32'd1;
     memory[11496] = 32'd1;
     memory[11497] = 32'd1;
     memory[11498] = 32'd1;
     memory[11499] = 32'd1;
     memory[11500] = 32'd0;
     memory[11501] = 32'd1;
     memory[11502] = 32'd1;
     memory[11503] = 32'd1;
     memory[11504] = 32'd0;
     memory[11505] = 32'd1;
     memory[11506] = 32'd0;
     memory[11507] = 32'd1;
     memory[11508] = 32'd1;
     memory[11509] = 32'd1;
     memory[11510] = 32'd1;
     memory[11511] = 32'd1;
     memory[11512] = 32'd0;
     memory[11513] = 32'd1;
     memory[11514] = 32'd1;
     memory[11515] = 32'd1;
     memory[11516] = 32'd0;
     memory[11517] = 32'd0;
     memory[11518] = 32'd1;
     memory[11519] = 32'd1;
     memory[11520] = 32'd0;
     memory[11521] = 32'd1;
     memory[11522] = 32'd1;
     memory[11523] = 32'd0;
     memory[11524] = 32'd0;
     memory[11525] = 32'd0;
     memory[11526] = 32'd0;
     memory[11527] = 32'd1;
     memory[11528] = 32'd1;
     memory[11529] = 32'd0;
     memory[11530] = 32'd1;
     memory[11531] = 32'd1;
     memory[11532] = 32'd0;
     memory[11533] = 32'd1;
     memory[11534] = 32'd1;
     memory[11535] = 32'd1;
     memory[11536] = 32'd0;
     memory[11537] = 32'd1;
     memory[11538] = 32'd1;
     memory[11539] = 32'd0;
     memory[11540] = 32'd0;
     memory[11541] = 32'd1;
     memory[11542] = 32'd0;
     memory[11543] = 32'd1;
     memory[11544] = 32'd1;
     memory[11545] = 32'd1;
     memory[11546] = 32'd1;
     memory[11547] = 32'd1;
     memory[11548] = 32'd1;
     memory[11549] = 32'd1;
     memory[11550] = 32'd1;
     memory[11551] = 32'd1;
     memory[11552] = 32'd1;
     memory[11553] = 32'd1;
     memory[11554] = 32'd1;
     memory[11555] = 32'd0;
     memory[11556] = 32'd1;
     memory[11557] = 32'd0;
     memory[11558] = 32'd0;
     memory[11559] = 32'd0;
     memory[11560] = 32'd0;
     memory[11561] = 32'd0;
     memory[11562] = 32'd1;
     memory[11563] = 32'd0;
     memory[11564] = 32'd1;
     memory[11565] = 32'd0;
     memory[11566] = 32'd1;
     memory[11567] = 32'd0;
     memory[11568] = 32'd0;
     memory[11569] = 32'd0;
     memory[11570] = 32'd0;
     memory[11571] = 32'd1;
     memory[11572] = 32'd0;
     memory[11573] = 32'd1;
     memory[11574] = 32'd0;
     memory[11575] = 32'd0;
     memory[11576] = 32'd1;
     memory[11577] = 32'd1;
     memory[11578] = 32'd1;
     memory[11579] = 32'd1;
     memory[11580] = 32'd0;
     memory[11581] = 32'd0;
     memory[11582] = 32'd0;
     memory[11583] = 32'd0;
     memory[11584] = 32'd1;
     memory[11585] = 32'd1;
     memory[11586] = 32'd0;
     memory[11587] = 32'd1;
     memory[11588] = 32'd0;
     memory[11589] = 32'd0;
     memory[11590] = 32'd0;
     memory[11591] = 32'd1;
     memory[11592] = 32'd0;
     memory[11593] = 32'd1;
     memory[11594] = 32'd0;
     memory[11595] = 32'd1;
     memory[11596] = 32'd1;
     memory[11597] = 32'd1;
     memory[11598] = 32'd0;
     memory[11599] = 32'd1;
     memory[11600] = 32'd0;
     memory[11601] = 32'd1;
     memory[11602] = 32'd0;
     memory[11603] = 32'd0;
     memory[11604] = 32'd1;
     memory[11605] = 32'd0;
     memory[11606] = 32'd1;
     memory[11607] = 32'd1;
     memory[11608] = 32'd0;
     memory[11609] = 32'd0;
     memory[11610] = 32'd0;
     memory[11611] = 32'd0;
     memory[11612] = 32'd1;
     memory[11613] = 32'd0;
     memory[11614] = 32'd0;
     memory[11615] = 32'd0;
     memory[11616] = 32'd1;
     memory[11617] = 32'd1;
     memory[11618] = 32'd1;
     memory[11619] = 32'd1;
     memory[11620] = 32'd1;
     memory[11621] = 32'd1;
     memory[11622] = 32'd0;
     memory[11623] = 32'd0;
     memory[11624] = 32'd1;
     memory[11625] = 32'd1;
     memory[11626] = 32'd0;
     memory[11627] = 32'd1;
     memory[11628] = 32'd0;
     memory[11629] = 32'd0;
     memory[11630] = 32'd0;
     memory[11631] = 32'd1;
     memory[11632] = 32'd1;
     memory[11633] = 32'd1;
     memory[11634] = 32'd1;
     memory[11635] = 32'd0;
     memory[11636] = 32'd0;
     memory[11637] = 32'd0;
     memory[11638] = 32'd1;
     memory[11639] = 32'd0;
     memory[11640] = 32'd1;
     memory[11641] = 32'd0;
     memory[11642] = 32'd1;
     memory[11643] = 32'd1;
     memory[11644] = 32'd1;
     memory[11645] = 32'd0;
     memory[11646] = 32'd0;
     memory[11647] = 32'd0;
     memory[11648] = 32'd1;
     memory[11649] = 32'd0;
     memory[11650] = 32'd0;
     memory[11651] = 32'd1;
     memory[11652] = 32'd0;
     memory[11653] = 32'd1;
     memory[11654] = 32'd0;
     memory[11655] = 32'd0;
     memory[11656] = 32'd1;
     memory[11657] = 32'd1;
     memory[11658] = 32'd0;
     memory[11659] = 32'd0;
     memory[11660] = 32'd0;
     memory[11661] = 32'd0;
     memory[11662] = 32'd1;
     memory[11663] = 32'd0;
     memory[11664] = 32'd1;
     memory[11665] = 32'd1;
     memory[11666] = 32'd1;
     memory[11667] = 32'd0;
     memory[11668] = 32'd1;
     memory[11669] = 32'd1;
     memory[11670] = 32'd1;
     memory[11671] = 32'd1;
     memory[11672] = 32'd0;
     memory[11673] = 32'd0;
     memory[11674] = 32'd0;
     memory[11675] = 32'd0;
     memory[11676] = 32'd0;
     memory[11677] = 32'd1;
     memory[11678] = 32'd1;
     memory[11679] = 32'd0;
     memory[11680] = 32'd1;
     memory[11681] = 32'd0;
     memory[11682] = 32'd0;
     memory[11683] = 32'd1;
     memory[11684] = 32'd0;
     memory[11685] = 32'd1;
     memory[11686] = 32'd1;
     memory[11687] = 32'd0;
     memory[11688] = 32'd1;
     memory[11689] = 32'd1;
     memory[11690] = 32'd1;
     memory[11691] = 32'd0;
     memory[11692] = 32'd1;
     memory[11693] = 32'd0;
     memory[11694] = 32'd1;
     memory[11695] = 32'd1;
     memory[11696] = 32'd1;
     memory[11697] = 32'd0;
     memory[11698] = 32'd1;
     memory[11699] = 32'd0;
     memory[11700] = 32'd0;
     memory[11701] = 32'd0;
     memory[11702] = 32'd1;
     memory[11703] = 32'd0;
     memory[11704] = 32'd1;
     memory[11705] = 32'd0;
     memory[11706] = 32'd0;
     memory[11707] = 32'd1;
     memory[11708] = 32'd0;
     memory[11709] = 32'd0;
     memory[11710] = 32'd1;
     memory[11711] = 32'd0;
     memory[11712] = 32'd1;
     memory[11713] = 32'd0;
     memory[11714] = 32'd1;
     memory[11715] = 32'd0;
     memory[11716] = 32'd1;
     memory[11717] = 32'd0;
     memory[11718] = 32'd1;
     memory[11719] = 32'd0;
     memory[11720] = 32'd1;
     memory[11721] = 32'd0;
     memory[11722] = 32'd1;
     memory[11723] = 32'd1;
     memory[11724] = 32'd0;
     memory[11725] = 32'd1;
     memory[11726] = 32'd1;
     memory[11727] = 32'd1;
     memory[11728] = 32'd0;
     memory[11729] = 32'd1;
     memory[11730] = 32'd1;
     memory[11731] = 32'd0;
     memory[11732] = 32'd1;
     memory[11733] = 32'd0;
     memory[11734] = 32'd0;
     memory[11735] = 32'd1;
     memory[11736] = 32'd1;
     memory[11737] = 32'd0;
     memory[11738] = 32'd1;
     memory[11739] = 32'd1;
     memory[11740] = 32'd0;
     memory[11741] = 32'd1;
     memory[11742] = 32'd1;
     memory[11743] = 32'd0;
     memory[11744] = 32'd0;
     memory[11745] = 32'd1;
     memory[11746] = 32'd0;
     memory[11747] = 32'd1;
     memory[11748] = 32'd1;
     memory[11749] = 32'd0;
     memory[11750] = 32'd0;
     memory[11751] = 32'd1;
     memory[11752] = 32'd0;
     memory[11753] = 32'd1;
     memory[11754] = 32'd0;
     memory[11755] = 32'd1;
     memory[11756] = 32'd0;
     memory[11757] = 32'd1;
     memory[11758] = 32'd1;
     memory[11759] = 32'd1;
     memory[11760] = 32'd0;
     memory[11761] = 32'd1;
     memory[11762] = 32'd1;
     memory[11763] = 32'd1;
     memory[11764] = 32'd0;
     memory[11765] = 32'd0;
     memory[11766] = 32'd0;
     memory[11767] = 32'd0;
     memory[11768] = 32'd0;
     memory[11769] = 32'd0;
     memory[11770] = 32'd0;
     memory[11771] = 32'd0;
     memory[11772] = 32'd1;
     memory[11773] = 32'd0;
     memory[11774] = 32'd0;
     memory[11775] = 32'd0;
     memory[11776] = 32'd0;
     memory[11777] = 32'd0;
     memory[11778] = 32'd1;
     memory[11779] = 32'd0;
     memory[11780] = 32'd0;
     memory[11781] = 32'd0;
     memory[11782] = 32'd1;
     memory[11783] = 32'd0;
     memory[11784] = 32'd1;
     memory[11785] = 32'd0;
     memory[11786] = 32'd0;
     memory[11787] = 32'd1;
     memory[11788] = 32'd1;
     memory[11789] = 32'd1;
     memory[11790] = 32'd1;
     memory[11791] = 32'd1;
     memory[11792] = 32'd0;
     memory[11793] = 32'd0;
     memory[11794] = 32'd0;
     memory[11795] = 32'd1;
     memory[11796] = 32'd0;
     memory[11797] = 32'd1;
     memory[11798] = 32'd1;
     memory[11799] = 32'd0;
     memory[11800] = 32'd0;
     memory[11801] = 32'd1;
     memory[11802] = 32'd1;
     memory[11803] = 32'd1;
     memory[11804] = 32'd0;
     memory[11805] = 32'd1;
     memory[11806] = 32'd1;
     memory[11807] = 32'd0;
     memory[11808] = 32'd1;
     memory[11809] = 32'd0;
     memory[11810] = 32'd1;
     memory[11811] = 32'd1;
     memory[11812] = 32'd1;
     memory[11813] = 32'd1;
     memory[11814] = 32'd1;
     memory[11815] = 32'd0;
     memory[11816] = 32'd0;
     memory[11817] = 32'd0;
     memory[11818] = 32'd1;
     memory[11819] = 32'd1;
     memory[11820] = 32'd1;
     memory[11821] = 32'd1;
     memory[11822] = 32'd1;
     memory[11823] = 32'd1;
     memory[11824] = 32'd0;
     memory[11825] = 32'd0;
     memory[11826] = 32'd0;
     memory[11827] = 32'd0;
     memory[11828] = 32'd1;
     memory[11829] = 32'd0;
     memory[11830] = 32'd0;
     memory[11831] = 32'd1;
     memory[11832] = 32'd0;
     memory[11833] = 32'd1;
     memory[11834] = 32'd1;
     memory[11835] = 32'd0;
     memory[11836] = 32'd0;
     memory[11837] = 32'd0;
     memory[11838] = 32'd0;
     memory[11839] = 32'd0;
     memory[11840] = 32'd0;
     memory[11841] = 32'd1;
     memory[11842] = 32'd0;
     memory[11843] = 32'd1;
     memory[11844] = 32'd1;
     memory[11845] = 32'd0;
     memory[11846] = 32'd0;
     memory[11847] = 32'd0;
     memory[11848] = 32'd0;
     memory[11849] = 32'd0;
     memory[11850] = 32'd0;
     memory[11851] = 32'd0;
     memory[11852] = 32'd1;
     memory[11853] = 32'd1;
     memory[11854] = 32'd0;
     memory[11855] = 32'd1;
     memory[11856] = 32'd1;
     memory[11857] = 32'd1;
     memory[11858] = 32'd1;
     memory[11859] = 32'd0;
     memory[11860] = 32'd1;
     memory[11861] = 32'd0;
     memory[11862] = 32'd0;
     memory[11863] = 32'd1;
     memory[11864] = 32'd1;
     memory[11865] = 32'd0;
     memory[11866] = 32'd1;
     memory[11867] = 32'd0;
     memory[11868] = 32'd0;
     memory[11869] = 32'd0;
     memory[11870] = 32'd1;
     memory[11871] = 32'd0;
     memory[11872] = 32'd0;
     memory[11873] = 32'd0;
     memory[11874] = 32'd0;
     memory[11875] = 32'd0;
     memory[11876] = 32'd0;
     memory[11877] = 32'd1;
     memory[11878] = 32'd1;
     memory[11879] = 32'd1;
     memory[11880] = 32'd0;
     memory[11881] = 32'd0;
     memory[11882] = 32'd1;
     memory[11883] = 32'd0;
     memory[11884] = 32'd0;
     memory[11885] = 32'd0;
     memory[11886] = 32'd1;
     memory[11887] = 32'd1;
     memory[11888] = 32'd0;
     memory[11889] = 32'd1;
     memory[11890] = 32'd1;
     memory[11891] = 32'd1;
     memory[11892] = 32'd1;
     memory[11893] = 32'd0;
     memory[11894] = 32'd1;
     memory[11895] = 32'd0;
     memory[11896] = 32'd1;
     memory[11897] = 32'd1;
     memory[11898] = 32'd1;
     memory[11899] = 32'd0;
     memory[11900] = 32'd0;
     memory[11901] = 32'd0;
     memory[11902] = 32'd1;
     memory[11903] = 32'd1;
     memory[11904] = 32'd0;
     memory[11905] = 32'd1;
     memory[11906] = 32'd0;
     memory[11907] = 32'd0;
     memory[11908] = 32'd1;
     memory[11909] = 32'd1;
     memory[11910] = 32'd0;
     memory[11911] = 32'd0;
     memory[11912] = 32'd0;
     memory[11913] = 32'd1;
     memory[11914] = 32'd0;
     memory[11915] = 32'd1;
     memory[11916] = 32'd0;
     memory[11917] = 32'd0;
     memory[11918] = 32'd1;
     memory[11919] = 32'd0;
     memory[11920] = 32'd0;
     memory[11921] = 32'd0;
     memory[11922] = 32'd0;
     memory[11923] = 32'd1;
     memory[11924] = 32'd1;
     memory[11925] = 32'd0;
     memory[11926] = 32'd0;
     memory[11927] = 32'd1;
     memory[11928] = 32'd0;
     memory[11929] = 32'd1;
     memory[11930] = 32'd1;
     memory[11931] = 32'd1;
     memory[11932] = 32'd1;
     memory[11933] = 32'd0;
     memory[11934] = 32'd1;
     memory[11935] = 32'd1;
     memory[11936] = 32'd1;
     memory[11937] = 32'd0;
     memory[11938] = 32'd1;
     memory[11939] = 32'd1;
     memory[11940] = 32'd1;
     memory[11941] = 32'd0;
     memory[11942] = 32'd0;
     memory[11943] = 32'd1;
     memory[11944] = 32'd0;
     memory[11945] = 32'd1;
     memory[11946] = 32'd0;
     memory[11947] = 32'd0;
     memory[11948] = 32'd1;
     memory[11949] = 32'd1;
     memory[11950] = 32'd0;
     memory[11951] = 32'd1;
     memory[11952] = 32'd1;
     memory[11953] = 32'd0;
     memory[11954] = 32'd0;
     memory[11955] = 32'd1;
     memory[11956] = 32'd0;
     memory[11957] = 32'd1;
     memory[11958] = 32'd1;
     memory[11959] = 32'd1;
     memory[11960] = 32'd1;
     memory[11961] = 32'd1;
     memory[11962] = 32'd1;
     memory[11963] = 32'd0;
     memory[11964] = 32'd1;
     memory[11965] = 32'd1;
     memory[11966] = 32'd0;
     memory[11967] = 32'd1;
     memory[11968] = 32'd0;
     memory[11969] = 32'd1;
     memory[11970] = 32'd1;
     memory[11971] = 32'd0;
     memory[11972] = 32'd0;
     memory[11973] = 32'd0;
     memory[11974] = 32'd1;
     memory[11975] = 32'd1;
     memory[11976] = 32'd0;
     memory[11977] = 32'd0;
     memory[11978] = 32'd1;
     memory[11979] = 32'd0;
     memory[11980] = 32'd1;
     memory[11981] = 32'd0;
     memory[11982] = 32'd1;
     memory[11983] = 32'd1;
     memory[11984] = 32'd1;
     memory[11985] = 32'd0;
     memory[11986] = 32'd0;
     memory[11987] = 32'd1;
     memory[11988] = 32'd0;
     memory[11989] = 32'd0;
     memory[11990] = 32'd0;
     memory[11991] = 32'd0;
     memory[11992] = 32'd0;
     memory[11993] = 32'd1;
     memory[11994] = 32'd1;
     memory[11995] = 32'd1;
     memory[11996] = 32'd1;
     memory[11997] = 32'd1;
     memory[11998] = 32'd1;
     memory[11999] = 32'd0;
     memory[12000] = 32'd1;
     memory[12001] = 32'd0;
     memory[12002] = 32'd1;
     memory[12003] = 32'd0;
     memory[12004] = 32'd0;
     memory[12005] = 32'd1;
     memory[12006] = 32'd0;
     memory[12007] = 32'd0;
     memory[12008] = 32'd0;
     memory[12009] = 32'd1;
     memory[12010] = 32'd0;
     memory[12011] = 32'd0;
     memory[12012] = 32'd0;
     memory[12013] = 32'd1;
     memory[12014] = 32'd0;
     memory[12015] = 32'd1;
     memory[12016] = 32'd1;
     memory[12017] = 32'd1;
     memory[12018] = 32'd1;
     memory[12019] = 32'd0;
     memory[12020] = 32'd0;
     memory[12021] = 32'd0;
     memory[12022] = 32'd0;
     memory[12023] = 32'd1;
     memory[12024] = 32'd0;
     memory[12025] = 32'd0;
     memory[12026] = 32'd0;
     memory[12027] = 32'd0;
     memory[12028] = 32'd0;
     memory[12029] = 32'd1;
     memory[12030] = 32'd0;
     memory[12031] = 32'd0;
     memory[12032] = 32'd1;
     memory[12033] = 32'd1;
     memory[12034] = 32'd1;
     memory[12035] = 32'd0;
     memory[12036] = 32'd1;
     memory[12037] = 32'd1;
     memory[12038] = 32'd0;
     memory[12039] = 32'd0;
     memory[12040] = 32'd0;
     memory[12041] = 32'd0;
     memory[12042] = 32'd1;
     memory[12043] = 32'd1;
     memory[12044] = 32'd0;
     memory[12045] = 32'd1;
     memory[12046] = 32'd0;
     memory[12047] = 32'd0;
     memory[12048] = 32'd1;
     memory[12049] = 32'd1;
     memory[12050] = 32'd1;
     memory[12051] = 32'd0;
     memory[12052] = 32'd1;
     memory[12053] = 32'd0;
     memory[12054] = 32'd1;
     memory[12055] = 32'd0;
     memory[12056] = 32'd0;
     memory[12057] = 32'd0;
     memory[12058] = 32'd1;
     memory[12059] = 32'd0;
     memory[12060] = 32'd0;
     memory[12061] = 32'd1;
     memory[12062] = 32'd1;
     memory[12063] = 32'd1;
     memory[12064] = 32'd0;
     memory[12065] = 32'd0;
     memory[12066] = 32'd0;
     memory[12067] = 32'd0;
     memory[12068] = 32'd0;
     memory[12069] = 32'd0;
     memory[12070] = 32'd1;
     memory[12071] = 32'd1;
     memory[12072] = 32'd0;
     memory[12073] = 32'd1;
     memory[12074] = 32'd1;
     memory[12075] = 32'd0;
     memory[12076] = 32'd0;
     memory[12077] = 32'd0;
     memory[12078] = 32'd0;
     memory[12079] = 32'd1;
     memory[12080] = 32'd0;
     memory[12081] = 32'd0;
     memory[12082] = 32'd1;
     memory[12083] = 32'd0;
     memory[12084] = 32'd0;
     memory[12085] = 32'd1;
     memory[12086] = 32'd0;
     memory[12087] = 32'd1;
     memory[12088] = 32'd1;
     memory[12089] = 32'd1;
     memory[12090] = 32'd0;
     memory[12091] = 32'd1;
     memory[12092] = 32'd1;
     memory[12093] = 32'd0;
     memory[12094] = 32'd1;
     memory[12095] = 32'd1;
     memory[12096] = 32'd1;
     memory[12097] = 32'd0;
     memory[12098] = 32'd1;
     memory[12099] = 32'd1;
     memory[12100] = 32'd1;
     memory[12101] = 32'd1;
     memory[12102] = 32'd0;
     memory[12103] = 32'd0;
     memory[12104] = 32'd1;
     memory[12105] = 32'd1;
     memory[12106] = 32'd0;
     memory[12107] = 32'd1;
     memory[12108] = 32'd0;
     memory[12109] = 32'd0;
     memory[12110] = 32'd1;
     memory[12111] = 32'd1;
     memory[12112] = 32'd0;
     memory[12113] = 32'd0;
     memory[12114] = 32'd0;
     memory[12115] = 32'd0;
     memory[12116] = 32'd1;
     memory[12117] = 32'd1;
     memory[12118] = 32'd1;
     memory[12119] = 32'd1;
     memory[12120] = 32'd0;
     memory[12121] = 32'd0;
     memory[12122] = 32'd1;
     memory[12123] = 32'd0;
     memory[12124] = 32'd0;
     memory[12125] = 32'd0;
     memory[12126] = 32'd0;
     memory[12127] = 32'd1;
     memory[12128] = 32'd1;
     memory[12129] = 32'd0;
     memory[12130] = 32'd0;
     memory[12131] = 32'd0;
     memory[12132] = 32'd1;
     memory[12133] = 32'd0;
     memory[12134] = 32'd0;
     memory[12135] = 32'd0;
     memory[12136] = 32'd1;
     memory[12137] = 32'd1;
     memory[12138] = 32'd0;
     memory[12139] = 32'd0;
     memory[12140] = 32'd1;
     memory[12141] = 32'd1;
     memory[12142] = 32'd1;
     memory[12143] = 32'd1;
     memory[12144] = 32'd0;
     memory[12145] = 32'd1;
     memory[12146] = 32'd0;
     memory[12147] = 32'd1;
     memory[12148] = 32'd1;
     memory[12149] = 32'd1;
     memory[12150] = 32'd0;
     memory[12151] = 32'd0;
     memory[12152] = 32'd1;
     memory[12153] = 32'd0;
     memory[12154] = 32'd0;
     memory[12155] = 32'd1;
     memory[12156] = 32'd1;
     memory[12157] = 32'd0;
     memory[12158] = 32'd1;
     memory[12159] = 32'd0;
     memory[12160] = 32'd1;
     memory[12161] = 32'd1;
     memory[12162] = 32'd0;
     memory[12163] = 32'd1;
     memory[12164] = 32'd0;
     memory[12165] = 32'd0;
     memory[12166] = 32'd1;
     memory[12167] = 32'd0;
     memory[12168] = 32'd0;
     memory[12169] = 32'd1;
     memory[12170] = 32'd0;
     memory[12171] = 32'd0;
     memory[12172] = 32'd0;
     memory[12173] = 32'd0;
     memory[12174] = 32'd1;
     memory[12175] = 32'd0;
     memory[12176] = 32'd1;
     memory[12177] = 32'd1;
     memory[12178] = 32'd1;
     memory[12179] = 32'd0;
     memory[12180] = 32'd0;
     memory[12181] = 32'd1;
     memory[12182] = 32'd0;
     memory[12183] = 32'd1;
     memory[12184] = 32'd1;
     memory[12185] = 32'd1;
     memory[12186] = 32'd1;
     memory[12187] = 32'd0;
     memory[12188] = 32'd1;
     memory[12189] = 32'd1;
     memory[12190] = 32'd1;
     memory[12191] = 32'd0;
     memory[12192] = 32'd0;
     memory[12193] = 32'd0;
     memory[12194] = 32'd1;
     memory[12195] = 32'd0;
     memory[12196] = 32'd1;
     memory[12197] = 32'd0;
     memory[12198] = 32'd1;
     memory[12199] = 32'd0;
     memory[12200] = 32'd1;
     memory[12201] = 32'd0;
     memory[12202] = 32'd0;
     memory[12203] = 32'd1;
     memory[12204] = 32'd0;
     memory[12205] = 32'd0;
     memory[12206] = 32'd0;
     memory[12207] = 32'd1;
     memory[12208] = 32'd1;
     memory[12209] = 32'd1;
     memory[12210] = 32'd1;
     memory[12211] = 32'd1;
     memory[12212] = 32'd1;
     memory[12213] = 32'd1;
     memory[12214] = 32'd0;
     memory[12215] = 32'd0;
     memory[12216] = 32'd0;
     memory[12217] = 32'd1;
     memory[12218] = 32'd1;
     memory[12219] = 32'd1;
     memory[12220] = 32'd1;
     memory[12221] = 32'd1;
     memory[12222] = 32'd1;
     memory[12223] = 32'd0;
     memory[12224] = 32'd1;
     memory[12225] = 32'd0;
     memory[12226] = 32'd0;
     memory[12227] = 32'd0;
     memory[12228] = 32'd0;
     memory[12229] = 32'd0;
     memory[12230] = 32'd1;
     memory[12231] = 32'd1;
     memory[12232] = 32'd0;
     memory[12233] = 32'd0;
     memory[12234] = 32'd1;
     memory[12235] = 32'd1;
     memory[12236] = 32'd0;
     memory[12237] = 32'd0;
     memory[12238] = 32'd1;
     memory[12239] = 32'd0;
     memory[12240] = 32'd0;
     memory[12241] = 32'd0;
     memory[12242] = 32'd1;
     memory[12243] = 32'd1;
     memory[12244] = 32'd1;
     memory[12245] = 32'd0;
     memory[12246] = 32'd1;
     memory[12247] = 32'd0;
     memory[12248] = 32'd0;
     memory[12249] = 32'd0;
     memory[12250] = 32'd0;
     memory[12251] = 32'd1;
     memory[12252] = 32'd0;
     memory[12253] = 32'd1;
     memory[12254] = 32'd1;
     memory[12255] = 32'd1;
     memory[12256] = 32'd0;
     memory[12257] = 32'd0;
     memory[12258] = 32'd1;
     memory[12259] = 32'd0;
     memory[12260] = 32'd1;
     memory[12261] = 32'd0;
     memory[12262] = 32'd1;
     memory[12263] = 32'd1;
     memory[12264] = 32'd0;
     memory[12265] = 32'd1;
     memory[12266] = 32'd1;
     memory[12267] = 32'd0;
     memory[12268] = 32'd0;
     memory[12269] = 32'd0;
     memory[12270] = 32'd1;
     memory[12271] = 32'd0;
     memory[12272] = 32'd1;
     memory[12273] = 32'd0;
     memory[12274] = 32'd0;
     memory[12275] = 32'd0;
     memory[12276] = 32'd1;
     memory[12277] = 32'd0;
     memory[12278] = 32'd1;
     memory[12279] = 32'd0;
     memory[12280] = 32'd0;
     memory[12281] = 32'd1;
     memory[12282] = 32'd0;
     memory[12283] = 32'd0;
     memory[12284] = 32'd1;
     memory[12285] = 32'd1;
     memory[12286] = 32'd0;
     memory[12287] = 32'd1;
     memory[12288] = 32'd1;
     memory[12289] = 32'd0;
     memory[12290] = 32'd0;
     memory[12291] = 32'd0;
     memory[12292] = 32'd0;
     memory[12293] = 32'd0;

    end
    
	always @(posedge Clk) begin
        if (MemWrite == 1'b1) begin
            // memory[Address[11:2]] <= WriteData; // Modified for task3
            memory[Address[15:2]] <= WriteData;
        end
    end    
    
    always @(*) begin
        if (MemRead == 1'b1) begin
                // ReadData <= memory[Address[11:2]]; // Modified for task3
                ReadData <= memory[Address[15:2]];
        end
        else
                ReadData <= 32'h0;    
    end    
endmodule
